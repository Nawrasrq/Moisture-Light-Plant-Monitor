PK    {�X�l�@  �     cirkitFile.json�]��8�~�����$E�d���`gL��%Q�Ƹ�^YN2��˜gڢ�ؖ-�t��ι4w�d���u�E�8��;7��U�&�\��V����ѽ���v�S:=N瓦��V�����G��4<:�W���͛	���L%$S&%"O)і3�眻�e�L�	ݼ�19Ñs �#NL���g��$!�%�)-��\Yemn�����'��.1�ˁ��<ɨ-2�g�"DnHF�"�L�ͭ*�Q0��-ӧ�sP�Ӳ����a��/uP�Ó:�|xR�s����'��G�LX�S�p+��@�h�`��0-3��D�O���9C�@�K$=�L@G�4�\Pb��Q:Mt�'�IGMVR!������L�`gs"
*H�ٌ�Т��:�g@�{h����E	m	�$�F�T�(�,�-��)��ɖ1ME�K"��$B�`�a6-yi�,-�i��l����#'GN6��l9�8��p��7�h��d�&���C4=�M�!hc���AMu:��u:�Bc:=�Lʍp�C���N����o:pn�}�,��լ���8�oh��H#X.|Ņ��DpI��"�p���q|�K���qYBWBF�h�3�\����2�Q�bC.<
���]��0�2�,i.*
}�2����g@p�q�������/;i6���l�@��NuR$���"+R�Ņ.4���A1�d�㠘�A1��b�<�yK�u6&�׍���$�C��v"4�=>�C��㲄���MVhz��IYB�����m�l��Ec�M��n��v�L��\x.I."
y�Kp2��rRG���Q.�����'cx.'Q��ṜD]p2�碢p�Q��8���8�eq������0��`�,�Y�8(�qP�#��8(�qP�㠘�A1��b�<�y'qP��Dqp2��rR��d��t���Ṝ�%8�sٕ����Ь��&���膳����v����殘@�VՅ�G7o��>*�9h�I�ZL�0�@ˁԘ�3ڸ}L�%�X�N�Y��� O��eд)�N�M�$�0�����:�l����Y���Nm0&��j1�2D�cT�XC�͘gm]��n����8��ջ)
V$�G5��rȂ�IJ���&<y2�5>��.0��p�!l<����7�r焵�r#���#2N���7U�*Y~���Pǜ�g'O�� �le�la)�S�3��G81G��Y�8������6��}�k�P����΋�,�-��l��o|H�Kd�G�D�xT�K䏟8����� ��H<[���2��HW�����0�� Q��B�r� / r� ��
N،K-]D�����\�r�L_���g�HV�=�H��l$�ө�t-��ŨP�5@�a=��	�R� Ohقq>n��y���I�Z,C�
��!"X�B���	`_d����Xk>>�/��|d=�"�]�E��s>Apu�5x�ȒC���\W��f��� ty�� ���E���>!�.�S��*�/���=�����h	i9-�W�&��Gz��v��#�8�P�M_A�c�}0D�t��������B;|Mi@���0�I��ב"gqK���)$�����¦B�5%x��eX�2,~��H(� ����,��o!��C���0Ϛ�X�r���ca˱��X�r,l9ָ���P�yb��Ab�}���|�h�&[�.��������;Gaf.��Q�t���f�u��~��l��OԀ��gj!��^��|��G·6>i��w QȤn��~�=h�Y�V�5���|]�+3_����jT�&�<����)�����{
�)�����{��S$�CC��V| �}� ��p� "�+ �]�q0Y=�u:��T�7�5�����$w��0�@}���aR��zܝ�C��{v.���Κz'��Α������sᇮ��^�Q�Cϊz�.jMvk��xf37��Ђ�~v͕WġMl��aQ�.J�ĺH�u�<,��"~X�����"�.R�Ez]�7v6��lO�e5�M�W����R"x
P+�&�g))�B
IU	f���O~���_,����c��C����ȉXӖBE^��'� �sO[(��S%��q�Af���@*��\�j)��� �pDg*%�['m�s��)��3����n'\|o�}l?z]W��n�����G%񢩧��@��}��}�x��Ζ�W»��|
-���}����;`:�)��@��տN�l�6����i��M��|YڼY֮>��n����������Xz�	^*�d�j1m�/.{�0u-��G��H��3���8�ό�#4�Vj�G��a�/%Ks�m�Qɯ�/N� 4o�<_1
��ǣ
z=o�J�Q��|Z�3�V�ۄ�k9&\v�N��m߆��ڝ�}��ڶ~�6o�e1�6]���������N�_�V�^��%5팪��Z�<c����IA���D	�K���,�O�TB� t%b�誧��7 �GQ��U�^wJ��6�?lS¨�)�-�]*%�EI�Jo�br�Jm�R3P�+u:ff�ޘ�A�S	1�I.�Tf�I��F:�"Ż�U���⺷O�sXK��Z2��
�e������*�o,��@�TK��Vt����P�SM�����֣�>��T�aO�>@�T�� 3%�uӆ"�7�R�qY�
W�?޶��vts;Z����v4�M���4唧�j��U:��UF���PFj��m}��qV���K�0{��e����$M-�� �@�A/����&-�o��>�?�1c�X�s.$O3�L�o�^����u�Yk��
H�,�0	a<q�Ԍ4]up�r���,~�1���.�=��~:+v8�i��p�l�QT[I\Z�`�m�iw(��u]5��|�K	#f3I�S~@���%I��,�=\��U�+M�'i�2|2�rmF�V ��4VSE�[���v^8O�= |�>B���?�3��Fn��}W�,�UK�[���(�-y]�ͷEQ��b]�i�Ƃ�q9��p]O׬� ���N*E���P-qb�Hf�ѥJ�(!�S�p�B��$��$QE�4�} �,K�U�������\Zdi�X���� ��)]�rJO8�2%.KXɴʴ�����ގ�U��j�����������՟�|�]�Q-�Uɕ�}u�j7�j��z9�� ��������W�hVU�|�t�æv��6�����l%�7sy�B���Ә�G+��W���� �U=!���o~��0���W��y���?.��cՕAO�������rm�;��if� ��9Ɍ�IixN����J��X5h�",V�I�cս�Ӏ�%��넯����fdo-#�#�yq�\�J��k�m������zZ
���z�̵n���o���ة����_zM�K�+�����t':���m�����l�a���|,�%�	X_�TJTiS�_B��3�*x�0����6�������B�N�^E߾ ���������X�b�%���J��B1���bH�T+�2�3�cNQk�"��EdY��0���!-<��ldk��l3�H���-�+�w�VTK?���T��S�Q��מ��sO3-�������tl C���B����U3W�K���V�m�-����>�]�{�׼���W�������[�'�jۃ����|�\}���z���|�uw��)�����Z�T�� �+)�$f�&�
� Ა���B�:�6l4d+< �Jz8���Vs�[��h���f�a���7�`F�5n�OӮכ����U�σ[�`��Mha�ʦ�,i��ħ-�Es�Y@�~��Շ����o����t��SG6�wŋ͎���5��N����'_yX}�(d�m&������ưn^O��|��O����yq�Uء��Um߿�)��!�t��t޼��}���ۑ� |U��o�Xh�?�y�_�����������X�Ժ�t;�8A�<� г��ўU��4r�I!�.�+�dH�A�BQ�.�h"��F6qQAcA��8W��Z�*_�>=0��<EF2���p�b�0�5]�U �I ��=oLX�x�Бa���B	,�+���˟i��]�U�`  ���a����n��s#,�1Q���F8�7��j�:��׎�T9SA:;+Y�k��~�xg*���?���hSu~��:m"<\�+E�!�g��}ՠ0�@��:ߨ��a�!� lP�`�.�3`[}w}HP%�4�K�G*��b���Qa4�ݨ�����p���f`O�!�X�,���Z�	�Jح�x6匈��b��/�8��Kzc`-�m���a���3�}�h�l��۰ }�U��~{d:��*����v��x�.�7���';_�ً��e���·w�F��PK    {�X��U
a6  \6  /   images/0287c76a-3da1-471f-86e7-79c7d2df61ef.png\6�ɉPNG

   IHDR   d   �   ��]s   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  5�IDATx��]|TU��OK�=!t]:��모+�׾�kÂ�.�J�}����������6@z'tHH�}2������y�d2�LB����%ɛ7��{�=�63:�V�|�&�`�#���2Z�P)���H��*ň�R��H)�rX�)�lv�:h�Q��K�/�4��!�| �����#e�0�\�9XJ,N| ������3��Y�0c���R�И�:n��/�ץ�Ç�<.��!J"�3���"�Z)����	��MR^��!�I��Aط�$�C�ҤL�r4��$�r��x����
�.�KyQ��R

n�t�1�f#ܝ�@c�,t1#�"�7L�CL��`6k&���	�݉&���{0��I��l)���@ʳRl.�HK��
w��Ky���2p5iL0������Yq�7N~�BFBb"��hifT�7��܊=y�ظ���Ub���:s�.�Ș��T�T�˵�5��1�UIP��2�� �]�MY=���ӺᲓ�0�W�������1��hM`ɤG��ϵ�x��<�=R��,]���<$e������IPf�HyI��"pQ�H38�^���OC��&ohr�P\�(�`Ci���"EI�!HKAjl(�"d��~q�����X)�Y��l�U�I��Kt�:sn�R͇�0�U��0#S���"�4~���#���s���?F�F|���l*Ŧ�(*���f��e�jq�LpB`		Cj|F	~1*	�ODZ|�b�oO�_���W���ïg#��N"!���p���2YJ.�Ŕ��a���d���Ԥb�y=��C���l�J<�a>�P �����1&�
���fC��!���e��Ʉ
kr�#��#~� SX~1&S/����o��.��{^؁s\�c����)J9��1�/C|��]�a�Y�ʒ[�`�%}<�w�����}�t}�bpM�d%T!�bW�;��,�.��'�	77!1ܪ�=�W>���-�ŗ[�qƷq��x���*���_>c4&L����@�؛.Ra�i� �UIiˆ0z]�񠢣B�����h%8ſ}�x��=�����A�X�7	�mS+jr��5�����2UW��={Of�z �M_�e�zIo�I����QSk�*O�4$-ϑR������d�+��NJR�h'�<�?nߏ��ø�bE`���r	s�n���;n�c��*|����>\�����es�	S�]%)��˂�d����f�a#��]�m�%Cg���Z\4g�u�0��l$�7�.�&7c�e�O|5��X�	3���#c0�{����
���T��E6�r�4i�8%ڗ)�T�)R���(�/ұ�֡5Ef�����4e��	{`6::�����ì�5a;��b������S����n��h�*]�k���xI]F�]Cqm�:���[�I5E��4g�֑��3G*JKa
�g��zH~�P}0���G/!�@�=�5b�����\�	��	kMPꋸ��.���r�K��JIc�Fo)�'!w��2����Xz�P�78m�%C{��B�Zqm�ճ��n^?*��2�6��@�щ��:l+I����ǘ�߉K|�0'�_}l�(���#�`���%_>:V�%��;�p�����ēwS�w�� ߜiLZ/���b��tdH���a��w��xS4�TS�$C��U��47!̺��"ׁu�iȩ���H0,���G���ƕB�/�)_�[�796���#+�¶o��������o�)���޸h����9�>��n���wm��h��Gk�9��6��R�u)Q����%%)`c:�8��M.m��h4175vH�;����q�<qm�M�f���lN���a��65��C�1*��R���T���q�+�-���|��gd=b���1�����[�5�p��2��XL�������X��<��i1�O,^�k��E!:ܬ�М�D��+��J����/��#�I�Y�,��K:8�qc�Ƙc�:�zD�h�U�	'�����(x�|�ϩ	�<sSF�� �q]�@̐ћ��0Mi�r�2V��&'��D��Y��^����Μ/(p�*�헺>�����@\���Q����Q
W��[�� z�t��/��u��r�%���B��+���sz�@���`˾
=�!͗� /�䖷�HK��+�Fa�x!c�������i�d�x0�A���U.���l.i����bTƖ�t#p}.�J�0��[8zE���K�xu�}jJ���3��Gla�a&Ǘ�$��\1��K�`��8\*8�=G�[e��&���	�(5'����N�]|:���^܁Tqn8�;���M}Ҝ�g����kZk쩛����ɸ�m�%rq\��!Jϸ��44���c�춓0|�*�E�y�|�קf ̝�en��F���>w0�G͛���;�����Q���E�;o%���!|3붘o�*W�)ĉ�G2�	I�>�`U�y����4k�'�D��ZLH�� ^����,u�n-|��IRJob���~�b���c�)�����_yP5HU5B��-��yb��5������N���{+�M�n������L^ݯ `�D��.q�;�b�d3txh��Ia�wl�;Ս���Wv��w��Y��Ǣ�ʸ������g�|���B���E+�$x��A�)mP����}E��M�l񭈴'���$`OD�'������Bd!.G��A����1���ԄP��7�k�	����D�r[���H�R�)_UUOo��!�f;��X�΂�")K��eR�0fn��5YTW��;ĉ�9v��t����P��Hg�V��0����a�c�����ɟǫ眵���JcL����o���?�k4k�b�rN�^h�P�d�J%�=<���q��^y]$<�S-2Rh�८������}����*���g̅P�%�Y�~���#�[��nq`bF��Z��=�U�I	s_č8W2����ZW[�1ۄ���ݒv���/F����,p&T��G����"��+eP�V�	�����9-�K$"93
�I��_��ή�a¯N�$� '}���Q}��O�pv� <*����CF���}�0�o�#����`�t��������#q%�t]ه�p�պ���~�f
8���,�gK��g}�F�с�(�����߇��7'��������RU�bc�>�;�m�O����xY�� �+������Au�#r����d^'�����`�����qXbt��j�b��u���'y�
�t�t�l3@4�B�&���`Q_N�h�NE��=%+\}��l�I]}V&*E*��n�_�FÌ��p�}��W����.���$�KO�"st�͊�0�_���{/�}��_��ݥ3�U����%����˾���k�Y�D܈#q%�dHzB��	�ϰ3�=��$g�8�%��0�^��Wv㥏��Be�&C����sMb#����r���g>8��?=��Ա���tE�R�nL�E�UVc��e�����#�a^!�UW�D�X_��6s�}N�ky�6C�>��w?�M���O+�j�˻�;�F$��,֢mV.�_�`()�+��Qb��'�c����_D���-Q��ӻṏ��Ʀ!`�k�64:Ղ1�~B1�U�*C��@��-�	Csl�q$��6�]d,���_ч��ث�j��y#���ͽ�˦�)�^dHr{:�O\Y��a@��H<v� ��m*��E�`м�@ѹ^}���6����ۚ;��������DkP�/�qz��sX�vd��ɐht�=�b��W���ս�-Rb����E'�H	f1�	a�jH��mٜ�)��8W�L��hkj�X�g�(����ś��ۛ��&C:����A��@U�����-�H���nB�{�H����ۗa����j�m���SS{��C�H\�b4��>42�#�h���}���؏I`{ �	j��ц���h�q�(�N��<q�G����GyC(R#<�w<��?1-=��(����x����G�;�\�%����Tgđ����n�'��@ix�����뱷�®R�f�1��������ke	9E:=�ޑ�I�3��dQ��!��#�Q�\Ѣf`CM��&����-?�,Ȓ�%���S�e}9�H�+q&�c���AiP*���!΋C%]���ʼQ��^L�6>y���s�")���6�à�st��5kcqa��pu^���d����xrN箵`�U6;zDW���7�Mc��4��y�md��ƀ'i�Bp��}����zj_o+���Sږ�����_ۭ�W ~h���QR�xL���ARgu(y�h	�>K@�-D�|D���F�I��ߐ��|w�wL�Zz�_5Vb��|?�t���	�;Zs@�;��rv� %$A��ݗ�բu?@V�5a�� �����W�M�E�&�_@�Р'i�Ƀ�-�V�0q��@��!�8sh�b���$3[$��&��xtlj�/��펅��̙���H�]>�{.��������Eܢ�3�jڌ��m��������
Ґ1�ʢ���ku�U��r5 ��/�o�����^*o���/P�����Ű�X]�i��S2��7�߭�o{2�/��0��ƧV�g`���mN۶�#�<���8�.��y���8����tL>#C�JX�C�p�6�1�ARў�9@_�Q�7�(_ۍ�ē�p��=p�����*q�3[�
�f�I�؊���N�~q���A��G0$��ﬡ��'�Ӿ���(KT�{F%��ͭ�¸�"H����.��;K�ߘ�p$0o�bu~�yHw��Ӫ���B�WԷs/]�ѷ�%%��ʉ�增�[����-gݿQ���T���74^G��T�H���Q�rfO���'V���"H�:��6���C����p�*���
�sT˂l����46�'I�o��i�����^
7�H �Ľ-� þ�Y���_��Gzr8*k�h�oj�n��Bb�̊�.艫��D� ��b���ݸ`T
��Ʀe*�qaʓ+�ڳ��%1s�����#Ÿ��Q4���"E
���?}�����.$�[���q�:Kx`�ē�[�Z[�2���X��L���!��L����P&�=n�N�̺,ekE�F���_��>i�j���Ww��/r�^Q�ۛ,��7�'��Ȝ��jb��0��&�גn��w��=��쇇0�~jZx��p��U�X-n��$���˞�s��azdʀ=_z���X4M�cR�taf��RLUJ�\�o?>?��<y�a�i�p㻇��oe�ǲ;)�ĕ8�XNJ:��rk���e�����Gbۡjl� �%!�E��[�����xw�E*~O��~���<��0����������U�����x��-�
�\�(��4���+a�w��rq�W��B���-���^#`rD~���s�2�g�:�9%��tzk��O��>�~~sV��������Ş1*+|��M�,i��ʑI��#��M-�h����^1Ό-�p�������+�c�u����b�W7��^�{+I1��J���e����S�D�p�P�]P����1~����)jy�0�dr�&��&qD��ʸ<�{L�-46-���D��ڢ��;/�hh2K�CЯO��nG��=m�hql8�g�onR��pQ���#H��5(�a�؉�e�q�hl
n:�'����c��'�C�B�$N@�H�\W�ٯ����+{��C�q�C,\�3v�J���IGj�S��C�j�������2P��VMč8ڹ�]�RLe���.�C��MZ9m"����oe�M-�_�e�ZZ���"9S��}⑜6�{UXox�,x{z�F�؅�����3�O߇`���W�ԸJct&0q�<���X<�agea������~|Xᆐ�oC���*hp/��z�bw?½ۗ&�����cg����ѳ7�ok���qְD��?����E)�>�M!y�x^$�r�_"�ا����z�Ig� �<(�j�`�!ޜ+�u�?����d�[�x�(�&N��rG���B:f|w=w�R��9%6v�!�NY%�Mq'���A�x�'1(�Aj���m�����Vv����S��[�բwo���"̋S��}��^��GSqŀ��Z��R|G;%�y+n�h��`�����x}� ���{\-3�/�N��&�|�*\��&�ƣ��DO'��{*��v4��!��Δ;�݊����8XF�SN��y#�D��o��aŞB�٣ #�ʐ,q	�O{O	plj�?����0l.LĪ�tXMi��E�0��>e��+e�|o����|��܊7>;���Ǔ~�jPLf>��>�Z�߭'�5�$�7�ݗ��K_��o��5�H�@��J	��a��Ѯ4��@�͂��P���ފ8�4ƣGZn�27��)1Ʊ-[$^�}�v��Z�"��Ѿ���8Cz�r�xp�L�N���]�W1%S�M�T�-eX�]�o�kP�� �Ҧ)o��K���/=
7���ߘ~1ʸ�PZmÒ�H~ ]�fa���`�t�9�6�l�"�y������አĩB`F��֎��&4��ꄇ+N|���A���e�I�3�N[r�0�pB1���}���v��.���+&f`�d$j*��=Kk�/z}��r��:�J [YѨ����:�p�A=�	U"o�����Q�ǅb��=<k`f4z���G[nш� �^E���j|�j���B"n�YN\F�p�2D%1n�RQc�bg~�R�}�ϼN�ї�z#�w�ae�'<C���^�����4v�K?�W1�<��<࿞!?7�CN0�CN0��3ĳ\� �����f��ci6`dV����ro�?0��YBΥ����1�_�щ�6��������N�><_<z
~
8����rCq���~ ������0k�9��k�Xf��7�'1���lm{���<��U���Vr}����Z��>r���p�pmm��Բ��9�!ɉS%�YS��qJa�ˀdG�f�[�HsS�ݳj��N�CFls���Ww���%bv4���Q�����ؤW��T�<�_�q�osq
��2B�i���d	���o���9u�U�6�E�:C>�\�g_��U�ߥ2_�O1D�u�S��-r Q8Ԋ��w�ҫ�ɈO�.8:��6�/<�W�s`�-¯z�2۹���¤K.��~lWU�M()< o)���ap�zնf+~7|'�E��g���,��uq(9���HIIi17�7�k6�`���o��7�2S���ɀ&����%%%hll����!��W�X�	���1Ύ7���M�m�T?�ы�p9���MB�S`4j��D�Z��+j@c�Q��l���
;j,HJ�+lTό&3��P��kc��m�DN�K)����������cGNĀ�"�M�����2�x4�V�\�ж��&�Z��s�q8o©�U��^!Iط�iÄT�	)&��<Xڂ���8��1�	�C{�+�\��L*����gX�F�ITy,:(������0�Q�F�K�z��E��㰉W�g.d����{�{��c�0�r�"����C�f��ƪ�Z���9n�~�Gg��:;���䵉�(�������\ԉ�"X,�v���Y�!�˖-��7ߌ5k���/FEE��{��	 			�2e��}	>|8V�Z�����!���������~�-6o�����?��w�q�.]���<�5��9�On�L���L��Gs������������=p�KI�a��0�(�Y�!<h�hlR{�]����O�a_��2�0��&��a|�Q�W��)qx%��N�1��V�8N�./��c���gŕ5�=��[x����	c�h�w����>�i�6�#�YҦ�I.�%�R|�f^�PW�C{�G|R�"���e$u�h���[J�ʇ���X��;J
�h�O;2H"�͊!F?��эKk�-r����#т�Y�ظ���X�}y�H=��HM�k�p��9θN�&N�����
'֫��Vp�h]JK�E�5`��R$G�����X��9ev��󂅠���-Zn(��wJlk���񘑙�:�r3��~��4��Q�]���~ϧE����Z G��)0�d�~�e�p\rF7̞4[�o},���<7���Ձ�o?	s~7P����x��ډ��q�z�7��ŬI#�����0�f�Pڄ��.��B0o�8%�i��[O��0�Y��(�jw�\�kh+K,���_91�I!j1w[��~���1�*�k�b�����Pm)��XB�;���{ṁ��Bo��F���z�s+7KG���)���-�O��%tT�S�*�;@F���\c��*|���1x���-碼�uB�r��:����i�l<n/�g��
e��y���Ko����3������;9M��S\�xB/7��a��+����놠��D2����K|�W(.��4ǞvNx�(Clw <҂�(�:����ƉuL���^�g�NXn�7�'�t13��);z1�	�u����Y���=��*����9x�ͽꂭ��c�|�h���fl�W���>Y��[!�{��a*����	x�l��ّ.�9��3M��?R\�'4C����`֕���>_m+Ug�<��E�q�3[�>��}c�!�.��?N�Z�����j�������E�Ex8�;��~��m =a��7������e��S��={*a��c����A�ʼx�,��p/m�l��}�󯶖"�PFnH�2D�)���8�4��6��0�3����t�K)������;�x,W��_l-Q6�'
�V7�^����<�	�|�0�1�g4������>���������#5A3��Q����:o�ٹї�}��� MM���["C2�p���j1�� ��V�q�����b�K���������79��͎2\�h���� 2��˴Y����˴���,�1<m��}p8��BT�Y�N�T�Zg����1T+��k
��ze�v�u�4���ڡ";&!�y^k���yJ�s���Mm�9q(�վ�Z��x���q$�݄9<�kMv��� #)\�q��C���	�]�t�-ޒS$6E�p�+ �?�ˢ._-�_����4+Gj'K5� ���Om�;2�>s&�� ��CEu�z�F%��^�^��Ҵ-kv�����]��}��A��S�A�zyW�����E�
̆1�c*K-���S׹�:-�KC�SX�Sg~�S'�gJ����@��w�դ��/�i-��^1���U*�5R��ҹE��0�;uw���Iۤ���^���uu�A�W���!.6.���<�35�^-��d/����95Ѱsv����P����SN��2!&Ҏ^1e�U��F�N�>����8�>� g
��FU��;E{�@H�-;zz�T#!̪f2yd`Q}WŢ�.R1�Ў��M�G�I)�8���T��%8+$���o�f�*�1�;�~s��4��y�È����w���i�28��$�#=Q(��[!��!�8(Ä�gũ��.����Bp c�W����h�h{�qL�Q���j�n��V���0����N��t���}e�B���W8��y}ⲾDl��@�er�9=r0N�]y�/>?�K�K�ĺd@�Oor�.��ju����wA&�4,�C��X�����1���*CȌDQKw�܌>"�l�����\�sx��/���f�b��ja2�������R�wx�U��Bu�T�Bf���ǍCw(��l���j�|�����(u�S2���H�u�^��y�@�W!��Ѻ��O�榚�ۮ�ͳ))Q_��Y{����9{�G�
��]��&8�ꟑ1T��.UȊ=�0�s��t����|��<���i?^�H��Lю4$-o��� x讀�;�������_f�Z�g�Ӗ���:1h�H������dt�ip_4Fi"S������V	D�ab�.�}�3��;��EB�/��J��1>�1ITŹ&�k���!:A�]ֱ�"ۋS�50�ݸ20���[MJ�5B����r����P{JD��B�B����d�]�@ZN���sH���$Cx�`�%%$D/��ib��#�ّ�o������U�Eԉ��v���H|;��Xa���U�O���ڛ�b�a@B�6ءl��{�Ja���7'�7�;��P���dg���jIC��I����~���%:�k�H��Վl��O���)b���
Q_�(�Tcܵ%��RpXb[%������^DZ�.4�A���b��R��E��Vo��h�&��p�6J�����xj����!�Y<�m��/E/����ȔSD���VJ�;���>20�U�t��[�~��ߣͽ|���[���,��������;��8��3����Q�� )�tD��@�}$��}���F�^�~��m����
�F�� !Ly��=ESҖ�5d��\.��"�hN�5�ɧ�>1M�ػ�}�YM�ۃ�g!�w�t`� �8?�$�H�$F0���x���[����.�[unsI
���Mnd�f?���%�;|W���>v�u���EA^|,8g�����B���"�<��3 �=���ɋ�E�L��䩿>5�7���wmIc?���9,e�7�
���Z~E*V������O�x5v����G�T&�L�;� �
�Dpy� ��	J��p��73txaރ���C�k�ml�%`������:YwP˸�}��*��^����� c���o�>c��;yO�����{�0i��E��r��)���X��S�� ��?U��
���2:6��:(�8I��#*(�|ń4�UZ�XG�Ũ���~��9s���;��.�	�=a�t��Z�6W>��ͷNH\�;&��ͻ�
�#��+�n����~�-i�S���d�ߧ����	"uUs������=�697��4��=H/K�H�{i��PI
�p�ô��*�4����NH�78�����wZ=��.�]�yRa��U�l$C6A3�;q}\L�"r	�w;�p 1%\1m,�|�����GLM��gj�z�'�� �g��Rۂ>qUhr�-��/�� ���*����[D��=m>�^r_��ϝ7S얕8$x�hd��e\W-e��f8 -�?�韔5�+�x_�-9]l�j��og,ě�f�E��UN�F�g	�zV\��@�e G�C��3Q�=����]�������&�|�6��=�TO�R/�l 1��_�yEFzD}��c���b��{��gR#�h��i<��}h�o����l)��)�/�3DDI�x�P�E�x<-A�y�Lt��n|Z>0M���9S��[jծ�h2�b�J�sd��!�������r�Ab�kπs"-�/��z���-T(��F�*{�������F�R8H�A�r��{����y�D�S�E-҉��s���i�1�[�T5��H�C7�񰁒�hEcZ�.]?�2['��̖�dM����J�Ώm�Z,���#�z`>�~���6��0��n�H��Uo�7�05ϋ�l�,�n��|	�tc��gv>-�<]<���$z��A��$Iu~Lz!.�Key�h'
Ӟ�U�>2Yg����8�	�5��J{����H�?<��n�������δ��J
�H�6����B�&mIc�A�����:)[����h&Δ &��zTQYw��鬴��Yא,�FˀJ5�2D�ׇ�Z��7�׮������%��!8pt�(M�H�h� U�,��XT�5�r�����d��O��F���w^�z}�!a����g�~����MRߛ��z�V�Ź �5��h�<�JkhX�ѹ�4��u��g`nu���R�5�B]["��Ǉz�������X�<q��F}+?��tR���Yî19/�n���+͢�_���,Q[��C:�{l׉*yY���r�M��_&�� ��x�y���.���A��K�O�ȀN�׉��f�5��B����H�^��Y��;Ȼ*zV�)i�30I{��ۅxC
]�$�O�BO��Aƛ)lH�R�iV�l�ۋ�F���1���vf{�~��h1̸^�	�<f�cD"�2�w1��~�[�ѽ��u�R:�9(�]��>L�A�!o��˔Y̚[��Z��zp@�)HW4����h�����2.YI�R�_�2SG�i���S����@��p���)���2E�9$��A�RZ�^�W{�����Kf�����w���#qۈ-*س�	�gPr@�����Ϝ̋R
ռϿ/uKȱϟ�r#�R�/��l��S،t�܌�|6���� �c�K?}�;.�h��.�}%#�sտ�ǓRq�97����	�ʰ�)�㜵T�*���u���-vM�f���g��H|O�U�fP:���VYiEJɤ��U�Y,tx����_��q����%*CCɕ6t��1��O���$OG|���s��W��E�2h�ʭ��۬���N�N��S�:!#_�ę���N�\63�k�3��hl�#��/�./��=a�6K��#��B{uw�b�/��H�b��Լ~K۵�Ms���CJ�o��� ���bQA����T[�S}�	pW�w�RQd�p]��sy�'1�
#ߑQ]"m������7��r�g�Ș����$D�H%���Y4��MT8��0������Zu��I�F}�����S�=��n��o��0��TN5�+��rlM�+���!�8S�.P�%x�ZsgA-����6�B�HK��q Y�0����x���$�:^5"�5��8���c]�X�$]:-$����_���/2z��dF_q_���0�O��9깘�����7����<:Á�]�"�|�O3�xI	��K<ie2:���)����o\%Ɖ��>�G��x����#3����RB�3��̣�z	��9�l���1�>�;~F��`n���e��2�c�,�ܗK�BJ:
�%O$��A���F�̕�N��🅽�h����_��$@�\)J��������t 3H�\�i�/�k���t�)�K�nt���9������U��?l��8#K;|�~T��/%m���'S�^��=��e��K��2��;M�������lF���5f�^lݜ)��JhIȹh�v�
��z'	��C�p�2:9����q�C����yƶ�An;Bs��!����Ta���%�ݽY*���ށ6o��͗w��?1PE1�[�a��(6㒠��a�n�1�$�4�S܍ϒ��	_B��DJ8�͹qfM��\�>���8o������6fp/'�9H�z��TxC����H��K�,�Ƙ��
c�x"����v�E}q�8L��L�W�L�s|߉d�ߠ1�P�f:���KZ�@D����WI�^�I_0��p�Ӱ� ��W�$��|U�?�1�a��u��j����n�:af0u�2IʹЖ�6[�g8�P�t�����
��n����08[����.�Ͻ$���S��xS�}$��P)���6.��B���`�ͳ:�p�����n �7Gۛ�XZ����K�/�?K4�'H���    IEND�B`�PK    {�Xyɜ��  �  /   images/110f4c69-ce42-4daf-8800-65b9db14e3fe.png�y�3���tQ����F���E'Z!����� !8D/�[⢝Nѻ��{��|g޿��wgv��}vv�_vgg6�P_�����DKS�:��� ��bJ*�����K�����������I:_5sߗ�N��0(F@@����[���^PAO�s��=c����q���W�AO�]{����s�|ǋ5���5$��/�}�6�av�B��0��Ѷ���*��� �mik��Tr���ArlIڥ�z�!��lS�I_������i�|�J��?��!�����"L�L�f�>M�8�~SP��v"p�_��b��*�i��:�����X*������#�F&~x������NG�2Jr3��?�P�sH�{�>7��<X�̠��A8po���k	l�ʸ�x�cu�����[o�Y|��r��q~>௳ .��P�m�^��H������e�/�����$��4i�80�o���j��C��ޒ�<�M0Н7!���[v\T���D��As  ����؎>��8;E*F�Z'�"�o��x+�G���Ǫ���8�i*7ls���Ef�;��&�f�o.)j(kX��㉉�4��`=M�¬�x�W��Z�Qj�5��.'%lNVi�����ZᏱZ>�O�.��鶭LP4�0��F�}�P{�����m�9��#e�I�NRۯї&G���k���ֈ�h�54�
��ܳ�=ӄNzۆI�<��ΰ �8�Ż&���B�/h�;ykm�|���ks�_T4�-:���Zt]:�U�QL��X�d�M�P"{L��<�8t=�º#�QR����{B�hh�-��j�>�
�V=��d����~�?}���Ԉ��˽���[PUS��H���,WkD |��k]��!��8ex�y!}:f� �TP�#�x��(�l��e.��9�.�G����qy���{�0�8�����y�VN� �t<x;:[_��E׫���O/(�����C ��/�D%��{�&���R�����Ȏ����l�	��q��9�g��0}�)���$+���<�����?��tl�3j�2�I'����ȭ�7�5zW��=��!HG=o�_��b-R������1ߧ?W�c?�&����l���'u��ٕi����QMrˏ�}�)8!�T�����_����������ƅ �fO����1���dG��
Y�jƁf�?
��"���F���3G����G��e�>2g-%�4����!�c��)��rB�Ƕ� �v��G��%G�a��PD�F�/�	̈́Xbz������?���-(�� O�vA��a�{�nq�iGᅂ�_�"m�j�$^�p!ZVgL���T������Nv[|�}NY��(�mFz�׃u�Ѝצ� >��,���svSBy�:�K����e���vx_�JX���k�|-�[��NZ$>����gR!;g��<��6�
���ei_(l�����9�LV3�֜2Q{�(�~[�蕇�Ld�"�gttE\ݞ���mS��bt;�f�&�P�c@NjB��aa~�y�&�����Q�X�
p���S�L�n\�f�3�E���s���'�쬨t�؛r�O�u�f�֩��	��t��:�Ȼ�V�����-��!:�	�P3Fo���I� ��cd 3�Q>��k54Kl�xg���sI�o	%������lJT�'����:�6Yd�7��e��|t-i"a9u��Z�������#�����_Y��W������P>�ɥ�פ}P�;�_)Tu����O;��Kw

%��,�%��yܔ����nH�ʇ=���Ҫ��p���O��,��Sf�F5��T��NOF��NKv22bh�p!q�ؓ�����I�%R�O��Mw��h;���i����Seͯ;� Hզ���Z��N��W�:iֱ��wy%�7q��>du)��b;a��3�y�0۞*�h�������`��V�}�0~��g�E��&�>�vR�_��=PΆ��W�4hiŦ�W��<�̿*�0��e��Vt����aG���.]Rdİ�p��b�]d����&O��U����@*��r��o��G���}~9͂T�.?�0�y��[�v�xc�>�sc�o;sӉa��1������6"?��[m���%�/��1�Xs:o��%a���2��D�w�~�S.Q[���?�=
�KE����� �$P�"j�8��v<~{dR�����j��l<1�T3�d��%~#�`>ߒ���IҙK�q�l�TS<֯x�po���\���׀l�ʡ��D���
R��A|2�jB<�τRX���� 1Rc��R,�mq���@Y1����ݞ/o�?a��c�2�.Q�t{�D�-k.C[������U��.D�,Z�3��Ge����x�\i�OWZ�	|�#�b�@��^���%�,_t8�|]���t-%�1�y��V�qC����T��žډx?�}Y�[>;*nn?ˌW��̡TO����fOM_l3�eg�K,WddW[�~Q�EZ�����FS��,c���g���ɭ	#�F�c�k���-3�����S!n���T��11v�՚�
�T�����O�480��X���S�]�`�X�RU�6ŘF�&^u�	J��1_)�@��$Ĕc�t�P�^$�%ETZ2�O��E�`�iN?$�֖f\Ծ��n�������Xd�hO����!�=�֊B� �>;�2������&M��4�J�
�4n���d)ЧO[����7]�$��tO28��@<FӦ�,&u�������DӺ��F��*?��#��ٌ�%f}ƚ����G�垛�@��pi(���L����@ӀT����5+�mA�ؗ��"t�RCR�o�1�n�Օ���A��_��ӵ���}i.(��M��`ܖ�	�ʦ�S��N�Ԩ��X@��r�ݨ�+|��mg��&'|�D�����l�LW�h�_ז�+&�`�C��gx�;�H��ӥ�v�~�L���k�x0j��8"��>�����;s��,	�w�ѫ9L�vE;��c���n-M�g�O�#�@�k�r�_�φ��1���w�/�~��N���S�f�u���X��[��N��%�DjK�r��9����� C�R��xtMM�Jfm#^��1/\�n�
�Η�jra�\h�1u�F=��O��9
�ʄ��h���~�>os�߫~�'Fw��D�����}\&eE�Ϳ
B%�ڰgF�F�j4���J7����s��sY3/����]��@)_r�T�Ǧ"�7��+`�R���dǚ�$[Tt�II{�\���Æ��n�n��q�^.�E0G���#��u���"z$1�p�а=��-Tf
�v$�&*VKN��Ɛׯg̋��ʹ�o��b�Y���������:K$��@t���P��E��h�+��,� ��P��z"5R�dEm�^�|����;�Io�G�&T�%7k�rĩs��^���j|!p۫��!�`Dn�f�%D'Ѹ����v�	w�� ��o��r�� FT
���7TTj;�@+	9��c�<ϟl��V�W*��U�����M�F���|o���6�b#���T��htl쮏�����2�`@9���<D�U���+o)�b�r��2pV������D^�O%��.�W]�����V�XDu#la���|k�Mr�����j�sG������P@�g�'#[�D��sWR tO�y���d��
�M�Ϗ��(���$+7�i���DmNß#_ah�o�~��h�c`8%���s��?�X�*���	�6�_~SxX�9>ZD(V�J�
�z�`6d!hN_�0�z_"*�� ��#�僖e��
󜳨���Q���C�k�'k�A�N�m8i�����QAW���V�ҷPH �@�\�Z�����v��a<�,A��T�I	h��߸V�87� �:M��N��͹Ji<|�kމ������sI̺��lE�����h,?�ܗ�Ӓ�m�?��t��a�!w�rJŀ�8��Kt�B�A䇋��x/�j�	L%kb}��/# _�7�օi�*[Z�� ���6����辧���������w�맛ʭ ���K11 G�M��G�2���O�Av���Ozy�8�l�\�z�Z~c4`&Tl���/Hs�^*�5xw��R�т���[Ű�n�-6�e�!�Y����z�a��NͰ�A��&��a��-���ZOR�;0�$n1��-��L��!^�)s��b�4�������Ϥ���`)�9z��k���8��⭍���
M��(��_}�ȅ�/OG;$�]����*>R��s
���1�ثq��(߬�SϿ��|���Q���<�T��dǡN�v���O�xQ���n�Y	cx_��utd������ϑ����|�#nd»�����b����r�Fs����J,�WV�v�������fs������f��n�{z���jꂕ�.񾾘Q"j
Z��d*4Sm"J9�[����>�zӜ2�]�R�S_�|��n�I7M$�{�(�M#��X�����]�T�ک��1�UP/t��&��^P3)�%Σ�~��~Y�.e�I���a���|��h�׉s�,� �̅{T!fg���|<����vC�4^y-����@���#1�1z&L�-ZH�<�x�TŽ�����#^h�����Ogs�;Ӫ�Ѷ}��f �CXmos��7�Jk� ��3u��r_�/gz����@�j��s6/�1��^~s�bٷ߿n1x�ɚH�c���$"����N��r�=�.�mYQ@f�lt,=��z��pm�(�x^�*�q�sG��<�Xϑ^zv'|4�+�[��-5����e[HaZ�E���)�*H1�LXpND~A%}�"�H�.u���]�����([��aT䝌�y,4q�@F�m!���<e �S>�=��c��Ml���p�p��~���Ώ�٧ѽA_���"�:'6h"7��]��>�����)�Y,��!x��E���2D�C |�3�������}3bFꢌ
Y]�p�qJh7gC�ʳL�2J��>2$Qk�7��*����V�݉5��	G\N)����p�rU�/��.,g��t��yM���n������Ȇ�
�kp��T(�MRS����+��jo�z'����"?4]��%��Y��N� �a�����}3İ���p�Nd��]�AH�fԋ��p���T�T�������C��Y��F��e�9Õ-a97�����|���ß�p��#n)y �d"uO��R��g�q��اv�_*�_��J/y�k��+�Y
���H��P��'ݞw%������զ<~qhzqzǋXÒ�j�R/�A�W�۔3�x����Wb#K&W����ښ��#L݌�ԛ1d:0�Ov����l'ں���s���g�eM���{4�?�'��Gڅ|P�%��s���T�_�V+�g�-��4�*�q-�8�{��s~l����R�jv\��y���;럘g��|�XZ���z����Cqfo��+�eG5��ځR���K>�m�Ic����_��P<����~�w}����B77�2&5�{���2SY�ONp��Yp�4����VI8Yd�T��Cq��I��1I�� ���ӭ����m 4�(�J3;Ml��o^� YMz����*~[�1���Y���b<o�wZ%�<Î�o�u�󪴩71��tsmO��$ٲ�U�8����\x�b�cWl<��T"T�����+R��"�]&i<���-a�ŮՕ��U��3���`�`�P��8�\
j6�����o���4���S�.�SƌK0���~��/q�>w
�q��I�@�7�y0=~��X�����i5=�%MI�P^���=��Za=�~�����dk`�Q^��$����ft2#/T��_���ihD�<�����y
[,�������T��o��sm2�b�#_^�l�ݞ���U���=���|���3�&���B�H���ľ���':���j�M�����~����k=�Ĝ�Xkt��������̈́��������a��K��On7�6�ӡZ��:s��D�=���������m�A�R3�{�Ղd@d��"����O�!|JY��6����(}�F՝����C�Q~�2j��z.06��A�o@�$^,������t'��Qw�X�^zY#s�;{t7�y�'��s��H��VʗlHEXJ4�-�O���jO�?P�_!Z�%[T!<z��VQ��.Y79��$��{�٤Ԩ�Ι��K�*�*̖pf^�,= �g^�^�f��̜U"3Ъti���Km�B+�?��8�����3�j*$˧��C�ϰ�y�]�����*�'d�V���h�v�2�h�uY�p���H�B/��Y?-^�i��uf�B�q���*��ƽ��e��Λ�j?�]��nD#�K���d�=�W�L4���1��������td�����3���0m5��XB�$KU*���>^$�֫�2�æ���U���+�߻}k۞���w�~ó�O���Yq٨摆M��|������/b��i����8jL�X�)��0S�;4��6����f��|�D����V��7�Y�؟�kk���&m=��� ���� ��2�T��J��fQ�Blՠg'ٜe?��|gF��%���eo�2�W�$y�^���U��n婎J�d����N���|M��D)4P }���F���u����M�=���� s�LN�#F<�\h.��fY��>/��6����%J�+w����"G:Ӣi����,�Aj5����IO�$P`�o�DZE�:��q%�W����W����bV� ?��m���C�@�f��@����4�Jr�^iSt:�Y�X\+�)�]�s7���&W'�!c�I��^�|>��`oْ�J�S�?NQ-��I|��b�]5.��b�l�D��Y��U�w|�_�D+vE}�u70e&�C�3u�&O��ڙ�1f����5�`Z	�)}������
�u8��io�(P��1{m_	\p��*X�RTX���U��i���z�m7�t�:�5mSy qR�����,n�J��3{�X�Do[��p��6�|�j�P�Z@�8�CpVKL�9@��|i��F�jL+$D�^�݈�0����j�^+�?��1
?Q��<����,]���c���V[��/�!%f����Di��;���o����V/{@O�����e�����:؜	�����Z���?PK    {�X�䓶� � /   images/132fbcdf-34e4-44dc-827d-09a965026955.png�wT�Y�/��QgPA�H�%PP�tA@zE�&]���E��@�H��~����ݵ~޻�]�����9g����}�9񉸡�u�����赫 G�#'/:�f`�(���5�C�:t�1����z���k �w������)?3?COG?�m�u�p����� ���JS:�@�E\��/�{i SB����[�?���s�?���s�?���s�?�����
c����A��?���s�?���s�?���s�?���s�?1..l������c����DQ�;1����9[%����-���w}��.'��3;�\�/|���Wh��ж�w���t�i�%��_��������~�j��w����P��S��OZB�v�3r�r��E�8:`7�h֤���`b�\�o��{"?���s�?���s���Fq�� t�t�k��iWg%��ZQ���X���9�G���N�Z����谥#�鏀7z7�;��]n[�PQ蚭0B⏣��/���t��/wetiD\B2�Z�QF�:�+auY��f\�@�;j����+������'F��~ӣ�+�qͪɱ����E$��@k�]�R���.#}��J׽��L:�Ʌ�?/ZE(W�A�*�>��,�gT��.���V��`/�Y6�l���g��G4��乄��6K�E�k5�	/��u��]TfTz�MDڝ�==����D��T��y���
��=���]��|�	e�i�f���k�N�O2"����2hە�,^�S�Y@�&���2zf��K���y�ۻm�ʵ ���sm���Ȅ�WT�J�=~�	Jqi���.��g���r�u�&����&�+
2"��u�����}�۫����<g��:��sB��?����
�m݁k֢�97�����F����KؑQZ��v��6?QTj�M��	thf*k��}H���C��ߦ������^0����hKR��AKC{�{|]9��3j{4��������Ur�t[Uǣsml��o߿l<���"Vi<H���xb�lr>%G'�+�`]�h�O��6�rq�3
�gbxN�\��il� 8�Kb�iՎez�����N�]{�Ҕ�-I��m-�dTy<,5PF�ɹ�hX�o���md�^���s{ç��~��~�,|��; a�i�7#��ċ�SB��:�.b�vUrs��Um�c�ٹn��I4/"�Y���l��0��&�U�ptY�MY9����T����v{�ڞ�}O|�H']�qA?�.#)~�J�.}�n���F�H��H����S�u�O�}�)u��Ӫ8a��{��%����;����m��k��SK���ɺ�sYw0�������,DsUz�l%�
��ʒ��q�G�1釠��``��m}��Zz����k)%i�򣰺��;�M�u�*�/W����z���I%1ԭ`�@��y��䪧�7�SmƮ�u����u[���\��G�Ud�ב�ڞxݎ�4l��M屵����{�w�h,�b���Zzc؝]��	�#����Q:)��	��^d��Gv7�����I!�q
��>������ƞ� ��`0�Z�-��%���F��ڒd=�,Rm��WvG�A
M?W����O��/�;����-U� �����x����ǲ�^ 7%b)޷R{:r]<��N_ ^�}a���� ����Xw��>Մ׌��2I΁/]X1"g�2���@΀�jU�ۄK�"�l��Urn4�&(�&���/V�����K�[�����7��>��D���B븹C&�/�٦(ԢO1jk����P7��Z���봵IN�����v�:I������mEZ5�=�3�b2�߃��g��p�����Hp?M:��9����v��;b��Qw�Rz�D�,c�J����wF5�z�sʪFW�}�ޢ2z���`�̬�J4Z�(�2�r<.�&��K \R���>u����is��U���O��J� ���Jޱ������!<o�KVI��\�9���/�1UF{Z���=-1"�)�H���h�P�F(�ȥ�L	lB�i�d�bՑЂ)��1����#��~r�����5s�/L*�$�}YI��l̵Q߀I�o�4�2>��IXjھ���x����p4��᲼���$$��7���i���s��\h�o���ڤDBC�ս�d�u��u"Q��4(�_#�U�4���˺��2O�s�A��V���ᗛ݇#d��+l3���pC��̮sc2TE68�Iq�BD_@e�Y��I����-�@�H/��
s��7�~1]��s%��d23�)ol�v�֏��)"f�l�o��3��������jD��Q~C�i#��#�Z�4���������F0�G�1cط��6����VeX�;��>��>fy��Z�v���|¹���7�d����#�
��d=�2��~ߵ�Ξ��L�U��5���O�����ۇ+���#v-�TM�/L�&�V��ѥ�޷tB���[�mh�9��V���D����\��|D��v�X'~�1�πY ���)����� ]q?�Ӕ�����<�6)�xz������Z��UlQHG�y�j���� �G �IH�/�
��5�@��b"M/y����7M���a}<g�VY=7_7�`���&�b>`��e�P~�Cy�lm.]}��K]�}6Pt�V��"#筬vr�;�\���T�UȜ�� ��C;H���T���r઴fQ�js��&�V��y�e�-�G�`d�H�l��8
N-ib�����pK���S�Sݳ<y��mo�u�� �LN����2m�d��4�WR�w�<�azcc+���gz���u������V�e����.9xy��u��A-�&?U�U��j{(r�D^Nx���f�7�$���u�LȠ.�~㘱���ҽ<�Cg���'B�^Zz�;�=���S���E�U�A�O��*�Jn��<��a�?�ܐ? 㿯�V0��kq=:Sr95���h��-nԘ>^6����:�J���4G�����%�u<���
Y'�=޳F�u:�z���%���U)[�/�{�*���V|��>�4�e3Rrx�K������j1| TDH��dx�+XfP*3M�,X (�`+�2$ X�f+��pE�zf �������Z 6�xx)������A|�[JUN]�.?ʯ�3�>쏣ו<�p�v?;�c�dI��U�Cbg�L�����1�Q��3;��]�+�_�],`�;ژ�Ņ)pu"�E{P���j���5~4��GѿC�A=:r�q�t7dwz���{�E�ȸ����<��_-�Лo��׏%�4��8mD���>��{%�ш$Id�[�eYk0�m猧d;�t;B*��>[y�-��rD��[�ab:˟�ܨ��|�x#pu7������}��m��=�5�Y�
���|f��5<�YL�L��TbA������u���E�I�U�A�9��w�SlM�3wI�����L��������S��qU�ɞ��ۛ�x�L0O��T����}j#)ֽ�`�:N�ҵ(��\5��Y��um�=�"�I��J�|ro.{�"4�
rI}�����ux�Ln���[�q��g���/�u��\I��ғVY�Q���K�!w�2�yre\X��'���B�*d����"����ȼ�*!F�AΨ�8�B��鹻z�G�M;萉_���!��OL�������}��3���)0�Γ+gA<5����%�X=b��C��`��лk��=���[c��{��އ�X����f\O����~�Q�����0aru�*�f� N$�\.[zh�p�5��˫�E�Q��
�t�Ū�p�o���s�q�~��5N]{�Ŋx���b�ߢ�y��<��dԣ�j�_�G�������a�R�}�$c���5gD����������#;{�;���a�R\�o蕱��9����)�BBҏ$+���D�1�!�ĝ�8��T�1��|�Y+x3
��65���o@<\��,�0U�a�kJȔ��?�u���XTG�N��{m��
0ZH����U�6�Y�պ���&����b�&��\����y�y5����e"N2gK� k��0�xPҩ�/��]k�WYn�]��@m�E�^]ꍪ�~�Y�frF鄩�p��0&�;��{��ڸ����W8���6�R���bb�:�P�#6U��ms$A(N�o�6(nU���[{��&�<{�pV�3��W��$A�:' �0G�L��Ě� ����<��U;�6����z�d1N�8������A�ʃr�;1��s��E$|rMu�7W�y��P=������O�X��q�Kυ�'-��#�{�x�$��c���=M�b��MP�Flv����������ݬ����`]���'�Ω�s�V+D�5T�v���^��f����j%m����f�� �A�|>Ӿ��L���d��L��v" ���r��,_�f�Z��?O|��j���]z�����<�������w�!������n#�05��lo���6Q�^ǿ\xsP��^�I�4��xc�UG�A3�O�dݹj%�/���`�������(����ҕE��v�}��*��s�m��`���wz�/'^�N�!�p65G�˝��Fj_��s�E��w��ǫ���Q`�*e�r�>L@��VE�A�θS.��&��P �]���LT�e�Y8��O�)�I������8[}��,�Q6�.���.t��.&e}//�l��"��]5�	ZSIE"F�����D̨r�N̎/2��I%�"4��+]���c�Sv|�(0�ۏ5�U�M�ߦ�x��q��4��C�,��uEQ�x�&�¿�$V�&ۖ(�0Q��)U^��Fa��4�Tgu+���sC��ͳČ$5�Y`dY�|���U.{���X0�1�1�>�2�/zi��xl�I�M��G��Mh �_�\VG�,�D3ކx���ƣ�0����ZI?�'��J������F��Ѷ������իn��A]�E�4��j go�\�H:93yBBT�7��Zn��Pha#1�>���L�j(�*x��ڌ'��+TEQҹ��Uв����{-��0���g�m�O@̖,T���mE,=5�C6�(b ĉ�E��
��L��T�R?��M��V�|3��I��M\�UПZ�iTF�1��1�1^�'h�CZGl{e�,�1��,���^�d8 �u�A�$����N�G�αCl�ɮ��Sv?����˙�g�A�NX4�]���o�!��쌢�wYA������&��V~�܍�Q��`JϏ�nG���=#�lf�ٴ¶c�`w�X��� ��x�ӥ�<A�KOC��x�@,��#�s�vO��!�c�(V���r>����}� \U�;��d������j˾x�^:nv�xN���i�Gb�n�p&=2�}�(.�!7�����[ ���W%��!��zr��D��!��lm��Z�rr<Q�?��B����#���o��+�[�nA�}!�7@��b�>~�/mR��쵫������s�y���_�`-8à>��q�V����q���2����g�r�n>|��f����Ĺ!�BB�cm�	3r��kiǞ�\$��e���/�.*�1`TغJ}u|�Qa@�y?�̛��Y���� 2�F��|O�"�C��BRa�׾6X�aF9�oV��B������Ч��	��4��<T���W.��Z"D��\y�������ƍ߇�i��#Jz;�!4���h�}��E9��I"��
G}x����<�E��g,�0���A��
��.�SE������
�A�l�}�6g��ةS�uk��>�ghi�=+������>��k��c��|�Y��1#n��8��&�N�<<Oj�CC+9�+K�WXᜱ���R���>A}�B�<k^�W�qW�4$���'P��B�a7�q·[�A2<�����VSѐ��z�B[�V2{sȢ���|�n!���p��)/&���ΑU�W���w�6��_u�E��]�\���O	����)�-���I�B�y�́_sԮF��)5_���9��ܢV��sͼ2��˖�U��U�>��dX?9S�����F *���'��:
lg!;눻����G�B�������W���쾿���H�sV�A�/�o�Q���MI�=����J!�tWl�U������F��&�y�A�NB:��%�Tf�#��5�-"�����^��_��z���@����!l�F�'�(�X�K�1*��ދ��dN=z�p}�$wE��G�n��+��- ��0	�=��2j�Z,*�-z`�	ic�hzf��R�����om��^�����Q��=��8F��$bxE5+H�#*i��1���7o,��޴��s�6��]�ƻ�Wn铲���U;� �e@��-�͌u���(���ֱK��v�LV,rQ�rGE�$[	��<�7�k����N�ċ�myxn�.r��/b�6
rm��h�{I��'����|���W��%��}N)X��o��P�z��X-�:�1}���{�����A�iH�	��km�{���t�M�^A�D��A
��QNb�DO��Q<2������~I�����g�7��P_�N���E��x>���@i1��~:J�BU>��K�\.�(�"��ē|e�^c���@�� dS������4�3�{�'�<k��=/�>$Z�AQ�-������GĨ����P(������=�$���9V�qp�,�y���o~�]�)=����	 �ziC���u�7����J�~�JUE\M�T��Dq*j�^ �~�N��T�5�L���O��1+K|[�x�s:�Dm�My;�W�����~;��	�zO�Ჺ����!�2�bc(Fq]�<b���v��*!#_�ַ�҈%��]P> �E3h�MT�
^8��ӳ�~�6g'�#\��\g#�7������v1��������\�<SG�_[ۏvx��J���d7���_� 4lご4��.$��l��Wn���OhŜ��[V���a��gM
t2���%S�ĬF�A� ��Bo�|�[�{GN��߾i�~��2�I��_�"Q�N��}���^&uf@�W����� d�"�i�,���z��ؙ9N톀,�`�mF������I����o��l�4Tx��W1�M���?Cn��W�7����;z���T�glŜtH�ߝ��'C�!��?TP��C���������"
)<۶�1���4����y�^�v�yw~�t�ze�f�5�{!�Aslgc-�Ge���@)�ϡ-��z��*��8R�����Q9��[�Q������L�K��W�%u��}18��v@ա�hg��}{{�GyF�Q�Ql���7pc>��Z?Z���������(�\�|��$���5������wh�G6pg1P��8�c�?'�u[=�J9{��L	��I�-���ݭ��?rk{��܃nھ�X����@P�p#���޳SB�&�ˤU8�ؒ�?`=���Z�$�8F�|�=�⋠���	-Y����у�^���}$�u�ۊyj��yx-�`�Q���Lp�Q\*��@��aЄ��t?���jp��DNj$�LqV3,9�R���O݆��;3q�(��5������n�x�b:�!$�a���26����(J總,�=
�0'�ϋ���!+�TRPPWJ/�>��T�L��m�~@���jnI�݅{�4&D��
��ܔ��4�������$À�"}��q(� TAG��4��K˪���p���A,�o�\j���|�D/?�3���y��@>`��L�9�K+��W��Դ虬87�ڑI3�a����$}��
E�,�
o۷xŊ}�@F�X$@E.\��rf���R*�1���x���>���\�L�����RSM�Q���yOX����C]DlvL�M�s;���cW�p(�ݞ>,Bw�^�?=��+��%d��}ˠW�Z��k��Qx�3� ��o$U\]���u��l'/�D����VP*q�`�k�Z�ݓ��V���i�D��C�N,GJ����)����4��Z�ɏ.\�2H�j��I�.�S��h��5��M����ʃ�A�)s���읔��_��q�uC��q�8w���.xm[)pm�bpm�I]�~=w0jZ�t��e���`���A��A��~T�>��j
$�mYМ4#p�?�#rg��'��Yh�;Hj�eWd��w���W
6�{Rs�[�`?�AMy�#:6�lyB��� q�ի��}_��6�=܉���j+)��� �L坏����j�)ۼ���3;��Y��I��7$o��������ZicD �l���ksv���VjP��l��&F���pd�&AM��m���-MG��*�̏��B��N�v��F�9�M�C�	�#�~2�����CsH��Q>3b�PڎSna*LY���;ڮۂ���H���"��O���#���/��K�Y���*��P�W>���k��m}iCkH0\r���	w�:��ua�3`��k�w1�`�~�M�U���ـ�}�!��;�`9����Pw^�X7�[�LU׶���v�cKѽ�a����!tf�NYL#Yv�	Du��#�y����̭�_mF�`���
����ka�ƥ�W��	��dj���T���ؤ\�[��\�W��]Q��תv���ci�wh�!�@Y�d�B��LU���5Ņq��Pw�Z�ж��^���a.�*%� �Z���rߑ�n�����_l�?��x�x������o��b��u4{Z���v�����αQ�T����WN��W�&���ɛ��I^۷Ѽ�Z������OT@]$��[��0��K5�@a���ۂ[ƀ�v�0K�F�Ԙ��Ǜ���˗�H��Ru��s��DH��/�DR���9�F��jS�A�&Md�f{U��f�M�B@;B���؄܌<5�/���:�+Bѳ�B͙�zaB(&Bf�F�#gԅO4��Ze�]{�n�eM9N�ʁ=U=�uKc@,#>�n�l�H:����f�Ǩq	4m��>�g���=��K�yG�^�~eM���1��Y�w����^��7x��V�&�����'#�8��=������rSQTQ�6hs�eʓ�\m�����gi�=֜~Ec_c+^!C�݄��?S1�""1����U��l"� ��/ w��6��Kk��1\.�����%� ��#�j�#72�C|'��l�����M�-w"������7�0�����h�#���>_cc�7+�����T<��0կp���l��^�6ȼ�:�r��|�m��x)����{U�;ӗÌ�Ƃ��vJ$��ڟFo"�¹�n��H�[��`��S�@;��$M���Y�V3�cY^�|�X2�w��wْ��;�p;F��jo}M,2x��FuǺ�w�@�=<��Su|j2��R�M_A����Y����$e�%�/9v�6\<9���8��@�m�tY��2̺� xmGvGi�L�J$W�[�����6���&���Q��Anv}�S�pb�8m{`rO��\:�N$�nT?����w�i	�n7�O1��"�;h;�΅~5�>jj�[įJ�(��J��e�/��}ȓ��=nAC����).�wd�V���,�\ś�������4D�p�vB��аo?̟k ~1M�&
65c��C\@��K�.�R�郹�,1�H�r`F��J�,�O�����G���U3wgiB�L�v�D��\"P/�6��%�f7Sm��+Ӝ)��|�g&��qKި"L�?��4���u��r�>T�lu�b�У��=���WoS���M_�F/��KH���җ�6$���(`��a%#$�Sc��[;t���9�~E\1q�b��'�0����@�e��|c#�i�+�]k}����j��s�h�W��&�@�v9|��J�֜��P�gZ���V1[�٬#'}�G���R��}��ؘ~5�mȚcJC�<����9������b�~~-*������2�5���K�*c�X�=Z�R��س���3�����^�Q��"J�o��sV�V�b�����dB�e��_��ձ��,P�ٝ�T����w�����kaJbm�ѱA]i���hK��ظI~y��G��&0$�!ɤ�X���9��d|@�Mu�3��0��%�@�Ѐ���X��a�	�&����N�we��M8k��~�<
�PYj;������?��t�ϱ(!�}�H�4 l��{�x���Y`�j�;�=��C�<��wd���&�{�n���POM%6�#��q�>�0#1#4���:��!�X�0U|+�Lo���A��3���Σ"��3=�t�z� _ꔭ�\�;���L��k�3{��d%��,����@p�U��}k����w� ��o.!��8��ɦw`Zh��wؗ���W:���}�^����z�?���@��MŁ�I^2���P<^�IcB9��������w�"_�S!'S�8�7�����P��
�EO��\��xbuݰ+��qߚ��;�<聲[�w�VS���{��� �N�f�@Ƨ��Eu��qb��T-ǴD�݁�$1����T3c��!�V_�:t���4�c؟�9`��ÖlObN=/�5g�>�U�6�Č�Ȼ[R�^f�� �.���0�{�=�(A��Q��k}{XkN1��X��`��NU��h��0Y�f���]=��y��5GoM������x�
.�t��F�v��.�F���� �e)z@��\�&��ʼ�}'7-qv�)������*�u(;չ*7gh�AM.E�!-��Q}Zި���e޳;�Y,�۴ẽ�֋����|�}{N"J�7��-u��T��iO����q�u�96c��{�|��
�N�AHk��m�^�T�X�'���x�����0�"�M�a=���Wvk����'�q�k����Q�:�C��.���nh��zu~��z�z��h: �-[C��6��N�ǻ��a�`�l�_Ā�q�:���2�i�F�Y�K:�Z��S�4�6�_E����&W�k]��z��I���g��׭��[�`�=T
l;�g���֓5���ꤍ��r����n���4vٛʦ&��*4c���q[:K��/�G滑8�7�M��=���'�m7�K�A&o�Lu�I�S�o�4���&���(�J�r6���W��o�?v��@��iWY���$�Wty^���eo�/U ���@����Q�ٞpG�{�/&&���=[4G��\p*�p��1l�A�A_��2y�3�/շ����r�޳���������l��.�\�V@/��	����?�/���_�R�#�����'s��]�x��[? M�[U,�'�3�u3��&c�ga׹�j� ?�+y;G��_oR xg+����՞	���Cg.*�󒇛�,�i�1Vr!P��Js�>��^]ҫ�؟�ZC�[:�z]>�R�,�<t?�K�`��Q�^r�]��]N�N\���&%v8&���I:5��aw��Ƽ����fڑ��N�q����=��zN�|C��g��c��?ί���@��s8��~_x�n����kJFy��Z�3^��6@��S��U@��_l�%���.�l�m�-�=�l�	8#9g�lX�۱9���D�9S*�:LDx��2&��c\
 ы���35b-��`�iA��l��F�Y�:��}P�ܧw�G���ge����y���0\��7\EG��e�*�CP�罟��N�<��z�k�uOLӝg�a�P	�+��;�r�xE{�}�F>�xQ����$C��%?��l�g�Li��X���)w♴`�ܩT��/F�)�@�<�����ש y��w����ea�a~����
(����Nb*���v)\�~E/	H�ŭz��?�Ԡ���^��}���������^D&7_���>z�-�� ol��8Oy����}-�[�djGY�� �9�M�'�-�~_��Ě^�U�z�}�o����9I�ᾈ&T=
���/7��*��"n�!]-Y���/$v��
ޯ����i�f�ݐr�^��!t��<��T���2�j^oQ_����u��߮]}'$�w}���j�\�@+n�7��$�VM��'2�!~@6R1��Ȍ�r��b=���f��J��ә#�$�K�-4ݒ(ޗ�}l��؇4�o@Y����߷ �����A �Q2�>��#e�[G~O���<R��!��n��*�케�$p���W_�2��zƌb躪Dj�1������]Z��G�J�eX8͕��U�Ž���M�a�ཡ� �p"�i�^Rm<!�T�S^^%g>qs6(�U�K�8�ӡ
A�~���^�p���o�I+�A�
D����8?EDM�d�"Ԗ&�V�Ӯ�I��a}����-L �M�������f$qx����):��"Fف��j����o�7���K����#EOJz�sC1����q�P]|�$�l-�bB�����#�gX�%d{X���m,��~cw#(^)謱�nMl>�@���yT�S�H"\�ˏz�S�VÇ��KaX�*�t��`䮘_B���>�X�Ȕ�ں�~0��t>.�
mj�6͎+��B� 6��n���bf	�Wkj��L��pZ���&�[�u���*���p�m3m:�-���q�D.�d6�;]W}'}�ϥ�Q�)E�۬X�j�>^�G��G˘�p�@�+�ڬ���(����ΰ8:O�J���ĖL�y�JC��N�!�T��xQ���u���[l�A��O�C�%j�<�=����B(�R��l7�
���`�uf���\ bH8L��������I�r-Mȉ�*RPw���]��:��~\\t���/�^��zD��ފ�e��0��-*����۟>����9z/^��!~N��i�E6�����'�S�U��=�z���{|�p%����U�OMvU@	[���!�$���Q��]�[�{��biU������+�`�)���k�v�7��u_ؽk>Q��~�%_*yl|��a�ca����TG�577}�����-h��k�+���Q�jq?VY5ഝ����3`+�d*,y���,�[y��nN<��J]D��)�U_���� �~`�NU&�s՚�F@�z���������qS�� o�e��yJ[�*Jo��5fgO=��H*"CwR���� =^L�c����	6�Lxu� ��|��R1�b��'B<k���M��&����)����	�	"PO��~ rPγ�nO%h���VI�okq@E�g�ԟ��U`��*���L�xp��
�"i���HiA�a�Z"�ئ�ę���O�cZ��cgp��h��Ls��LT�R�2��vnI_���ǈ�܏{�� O�ߨ���\����o�ꘝ>���.��8��Rw8sJ��kj.u�5�*/��\_a˂_�=�?o��$�YC���w��lC�B��R{8�[�\�K���E�*�w���7 /��U3ơ&����0x]3�e�,C*۵ek�B��X&Ǻ/2��c���![Ҙ�3@-+zاK�-�_�#�~��
�/�i��73������gp\ԙ#��:��yb����(,�
j�L���y����%�@	��@��ˎ���2��}��.���?�j�j�˸
�8.�ߙ�ژT�/�ߘ�<P�������ŻN��	�-A�t�}�<��i>��tP�L���Y�ʾ~�2.�7�{��
�E0�V=��=Ӫ���/#�b�t�K3�1���N��?`@����z�D���$Ѱc���� ������c=�Ы����׏<������<��Z���c�;�2��!���� �u�Z#�ef5/W�`�m�'M�;�#bU���2��p��ѥD#�`/w�����~�ꈘ�>K=O�ݷ&m<�j���u��n~�����\�zt mp|���`"����1}�D�+2�/�Z��l_X=%^l�Lv]�&�}Ï*\aFj��ǎx&m��0�@�Y�Ws������&A�>�1�Ui/qs��Wb��UQ�s9-����}��Qf@�:��B����lA���2��͌�y��m�5;�z�޷�.��������ahm�y?#W������!�3�����T	�q�ά����i�Lu�|�h�3�c���U���M�?O��̔	{
}C�zu�s��ۂ����Mm!}(
�������uD?����\�����s�˙��{�,���:�XШ�}g��@APVN0�����մ�E�����<��R��GV

R�V~l�ϱ?�^���O)����l�<��:�����uKĵ�'��`�$��dr)�.��FID]�zP���LНC��/�\���"(gv�ٮ�f�o�S��A�:]V��;TrkZ�~��A�@mq�@���i������m�Ⱦ��yfMN�{S�U�Zd����V�%��`^���Z�Ic'w�����<,��^L���9Lb��쎑����(&�U@��e�io�!]n�ȱ6�(Gw��X�!b�)ڦ�xTTۨB����K��l\�/Z�o�q�nW� �l������&�,>����2��U�(�M)���?��{��xY>Gt?�̠%x*<����,�(J�R��+��oL���+Ø��c��wo�|,p(3Y��y3S¹d캣�=+��1����D�_��+�W��� 	����8��$bhF�v���aoj�_���y�I��ҕQ�X?f����;� ��R׶��������'�4�	o��6Kܻ�q�\���_��	a�k��6
��a�ʳ
��v��!��k7XD�2�y��P�İ.}4H�\�&��ˏQ�(֔89U�~-sM����M�`�x���Eu�L c{l��Qg�)�v��?!<'�)���*R�q�� �dwIp~�Pn���X�%�8�e�-�4�4�����&-��h�1�]�� ��t�3�ke�=�.���ϗ�k����m���@M��H�m/1��T!���>��Ie����3����u.Ļ�n-f3�J�:�ʼ7��0���1�8��g��.�h���Ȃ1(��J�ŧ�c��PA�Qǲe'���IƶZ���j�52� A�������xO��L�[� TPM�6����.�Q�e�}��v<�S��
^?vN���������8H$�L+}kbJ�Bf7cX�B�\l�J�3�����ȷ��M�ۯ��T�~P��T�1Y� �zo:V�8���v�~p Cf�;�>Р׏���$���p���jJ�5����I/P�{v,���^??Z�*u� �2բ�j��.�"3F��<s��F�<%���<z
k�8@gnX���XF�X�*�!sZ�퉙0WO�@��_�-�[2O�[�^��=r�+�m5݉y�>�<[�NGm��Z���VOn�+�$�G҅ 4R�VD|Ջ��o��ʄ�H�!�}���x2
$�O]���b�t%��׻�����!S���yB;8��OGϘ�p�Z�97t�h�ŵ>���!�2,����_�i�B.��틳/=Z�(d?�H6f�&�9Z��vo[�hL;2j0���Sb�vS�N�FG��X&��v�C������ e�R���'`�BE�;L��x�7�	r���~A�������F���MJz�Ci���(�'�,�=y��SW�0l����ۓ�RLY|u	�8�Yh���nf[�X�ڦ��
1�
��sUd:����E	��<���<Q1E'eM����h���}O�;)X@\1p�4j���AQ(� �YG��91�z�����Ў�H��7됆�H�:4x�> �ɱ�ڄ<C�տ EP�)� K�s󔸩VZ�[�)�#r���T�pӟw͝�P��Q*�W�
�#��o�����b��]jo!�̬��
��w�)k�G*r$�2��J��ǏQ�`s��!�?����������r�A����;�UA���<ٞq�A�x#��V�n��r�<�͖�mWF�
�L3n&j����
��
���R%���:Ef��J��ÿ�5�O�ɂ�]�q�@qZ^�:FIFW?��u��ILvC��M�߽V��;�#<W����I�N�"�z���})L�d�∃���s`��9�E�X]�C ����ՄDk�T����z���~<����J��Ob
-z�9�K���>S�ٟW!����a�6�<p���P�Ds6.)@Ԧ�٪�p4r�3 /�u�$��ؽGf�t�>�ws)�x�L�fy�A����wF�oѸm���N�F��ɇr�AL̎e�(oW���$��hpB���p��<�H{�ѿ4`�}����.x�?���-�Kѫ�/�m��v݁�?�5�4��Xގ��&L)5zW�`ypD��5*���L��su����BP��R�<x"L �x'��t��t�ٟ��(c:^��l�3[�}��;��uz+���4�$4��d�<�"�j��m�Y*g�{�9���<�(�����!��+�>��|%��8�Lz�j�P~�����&�:����ڋ��ֈh��̑�@1�C��.�I+����,�M"̰qS� }�Rt��U�����/��X}�̭��]�Y����xө3s���R�s��_ؙ=_s{��ʎ{{�����k�ɷ�)5aW�VQn�@ӥK���/M�X^c�Ŏno�j% �����6h&�=�j��j?�V��*�+/��n]r&O'oT�>δ)��5}Գ��2�NW����o�[q������.ϩ����')����M�e�Dt���_W�<�	���?8u��(0��T�I(���ԙ
�!:u�[M1�ߐ-��L�8J�׌rX����O��ob���P8�W�c��B��Y�>�	���7��@Z�������ax����� 7��\�Ce@%I�+�?p E���H�ItcV��U�/-MD4齾3�G[B�t{^ ,4&��A]�:n����y1\��ÌߗT�2K a#��;��hĘ�H��xU3�NR]̀�]�2�_��6m����M7�忸	��n֔��K�^�UC���@bZ}���9끨��J %�qE� ��gpYm�[A�zq�7�v� lۏ��~{�GE�7-���F|���]�������:�X��	+B��uI�e������뛽Y�.�R;�g�|�<Eu������ e0���NdJ���K�,[t�~��Ij�O��*��;�ܷ���g��F~`��8���6G��3:%�?9�l�g?%����{���'���#��ב�SL�M�__��xkd�YFh�]�9n��}i*L:�Nղ����t;���VJ��\�`ݻ�`�D^G�$k}�5?=c�cn�2$w7n��?r�c쯍��JQ鯩��E���Q/�!��%�1rtS��I����\��EL�K��r���\Q1(q�cH]T�פM�c ��|�nU_�*���Q�1Ǟwԧ]V��.sS.㴳�＆�ɞ�p8+��dE�+ O�ʶu����=a�:�i���4�����^3�5����\݃��w��Źz�����m����h�D3K�D����fy7�?EY1�]Ev�9Z����h]&Bp�H�/�QK�HE{��^�\Q3I(����`��f�C�N��ޝ;Zɲ��Dc޶ڼ��Y*|D��@b�4a�l8uى�6��������T�Σ�����ڠfV�f���@�zMm�z�<hs]��o����b�\d?޸?�C�Ό�.�qJ����ͭ�H& \�]�q�T���?�����&�L�s;t�l�?�����m��
�[���۷6cc�=���fhv4��������z�x���|���)KR�$%�%YO�%	!�d�'Df�t(E���c���5�0ʞe�����n0����>�������C3���}]������z�/
I�2@�◭(ݎ�פQ�۽���*�ȿ���f|-��[�V��Wo�R�3I,�I\��J�8�|�5�Wa�Y+�J��]���[�T� &:YRH���`7��n��H[������h<�n1�u��!��&z�}�����,f�?��V�u��C4���)k���J��d�������.����^{��gǪ��6�=����s��G�Ro�H[�ͪ
p�r^��P���r ' ��[/�#��.ژ�s�uc�B���Ǔl�A�up�:�Ԍ� _�m�q�XU�C�Ҏ�(�}���ϩ�����fV�P�I��a�!BUՙ���@���
!��\ۓ�c�o�ܙ��.9m�=��^�D���c�j����� ��&u�w."�W=���&��d�\�f]����G��Y��0.������F?*��Sk��]�wECx�;>>�Ґ�;"1!ٛ����9�+�VD�k�XgZjA�/t���d$����z����j����O�4@�A\�����8�5�Ur����@�@
2l:�*��(D_���:
�I����������j@ ����Q0���X]��I�E%�ox���3�p��8�۠m@<o�bPq͓Rv��Ǉ�[�#�"HlH M<l<������=r]C�rt�����a�L!ߟk{NU�pΌ6<qq1կ�M��I�N��ay����΀RQʧLX��;����2���\��-w)�?��'U�K�?0Rs���C�~�0P��$Di�+��L�Ҿ�TlU�� ���󠫘�P�	�drI�4E�[_��X ���B�qV��w�h�91�^o��l�fS9���S������*��<@+�7����s����ty�̥�� c��Q������ٲ��^ԥ���"N�0�<��xrU��t�}�����7+9��S���C���:�C�EM�v$�(�ٖe*\�)0��Â�hYYY�c������ID�pY�@��*%�m���jӱ�z���u�!.��k�̏w�y7�u���J:C���#��������z����&���a��i��������wUJ�=��mӍJI�gfc+���h���D���$�ښ���c����0�vPo9/{��[�y?cx��!�������L��b�J����vC��������/�������1K�s�į`�qBE��d���i��s&{[4?'ޅ��!Ấ�ib�@�n�.�r�Z�c�Nr0���~�����m��UNPC-m���-�(��L>�M4Ց�G��,Fuj3���<K���͸C��}"�lc�zI�`���T/����Q������L��⥖�۽�$+9G��0��ǾZ�h16�D.=�jϔ�t��K��Ѯ����L6�3Wl��t#��{V�3��!-D9�������(̄�PAa)�����˯ɥ'W;{�dw�.h
|���ht��-oxK��������50PB0��r��>-�?/7b�]�	�h�Ȣ�c�Hv�G�O�ٗ�6���T���q�O�q~f@%=�fLdA��G�	�7K�U,9��̍�׽ �S����6�z���d����6˝�="gc����yLZ���[�}>��#�/V
n�]_i�����h�p���^ �[�%ĉ�/JsH����	JVɰ�s%�{~
��L���=H3�Eή�a2���X]�҈�O��:�z��M�8�X�����y�6dOv�}�h�K]a���� ����M�/�FR���Q�'pu��J��J��uDD��U$-/ծ�7��1s���;�B g��B������!���_���{6��P�v5^ۉ�Px�K,K�8���ؕ�����.�yn'��T��H���_�C���Z����*X�WH(s{�^�֛�֩���̊R��24��<����}�����E�c���;]2������j���p5yX��y��|G���j�0�(W��e)�SF� �tKj���h��7 ��*m�%�C$L?Eo����\RX��g� 6]05卝���5�߷΃�<=��󥫫��(��RW�;��J��B?4��1���K��L��I��!��cL��ǌv�7:d��ʨڛIo���^"�=��)!��{�5@O�p%ۚ����]��T�XI݋ʀ��/WG��IV�+t���[�: �<��F��5ݩ�v�?x�ִ���[cϔL�N1>�E�����x��|� ����S��ҷ�S(��eHQԪ]n��?g�����_$��ٗ�J���|�z�#W,#7��i�O����7&sY�)���ߴ��2o��kl�
�^��b��mպq�Q�S��]�:���/їL�&��
��vO��6ٺ��"���'퓸�����Ih�I����}������{��`���3��w��Xt�pＡ����J�8Y��浦��{/OJj��Z��鈌P��4�.��/������9�Ō	O��2�VP��5r�0�j��|��Gk�9���7g��9E���aD*����1�d��Ȱ<���H����Zީ���m@Eu��+�'S�vڣ�j� �/�ڔ�\Is��@)�t�A��+1������be��=s������+�j�m	H�]<�ut�.�������χr���+̭�Z��H���q{6�8�漣��n���)���V����с�i� Z���z�<ڽ��
�`lѩ��s_�=x�}��*" ��F�OhiZ!u�G�j������\?�\~?�(�$reЖ��)W�'Ⱥg���$�����4و�W6��;j���l�i�N�`M�N��+ks��93�ӹ��I��F�m�s��SF�'T�)�pk�f�$� �R�p�dc�<�t�*D�*#"��i��㼑�E4�N�`o;��	 $Zi��H�0�[z���q����ߚ������9�%1GҸ�밬TI�ҰR9��)쨧,�S��f���f�91>z�yiB��7���9O�w����]u"�/>i�c�G�Ba6Z��d�������.�������e���L��Wh6;G�U`us��g+c��YG��k���ƑS��,TOH;�%�)���e�F$�A�P7�oM�Rk*-���k�����
;��XDA{Z��Zx���3;���EJy�	T�����С��E�*���3��IV��ӡ{��>|�λر���h٭�:�z��Ӫܾ��V�G~�8@<��1ض��U�#K�a�hVK���9G3o��2�b�RW,0�1�B3sd��c$5��Q��@�W�n6�xy]�_��Nox�~d��3w��Ґ��T�����S�>T2#�P6F���{X�B>rH�h{�|����R�R����	8 �]�=k�W�DG#�-�/�>�@OK�E�x^$������I[aw��:�ph�C�	�w���8�Ì��D[���=ȩA����5��[S�2�P�c��-���}bɐ`��dXgSl�5,�aL�+<�(}	a�����x[P���!'��,Ÿ[M?P:��$�-ӂ$s �s���F�(��h'��cƯ�
�mW�= ި�1\�X�?Tk�)JE�u<i���ǌ5_�c9��cհ$��'t�}��>3�"o\TS�^�%�,IR��_�^y����)��s8q��F�/��i1辗:��È"��3[ߛGX�����xU���H������=�=�B�!G�hFҋY�qC�g�j+��S�A�R<C�%6]98�����熘�_�
P�`��o�S�_4;�;N�ũ.?>��-ͷk�����h��Dm��
*���s_����a���:Z:�$Q��Q�����Z�PaDF�>����5`w]0P���XV�U4&���mL.Hx�;~���X\"� bs��>!���a7�1����� E��:�S�6[� �?T�<�����*����[)��#�r��N4���=�D�J����`���4������YY�̡��ry�ķ�&`E>����k��˚���ƿ��I��؟�2��V*���t��Y�i�d��P�b^�L/����'�����f_ʕ���#�弲d�� ���ݪZ���8�_��:i���3F��1�ՙ��z>M񭄢H��L[���+�KoHeQZ�<𓻮x�'O_L%of��N�	n��~[)#��	���Y7
��k���3��T�*��]7����D�*���g��g-?�fl0�<�4�\VF.���]�M��HIp�B�>��Q�m@�'��rgAjd�m��(�,$XW���5C�!�l�>q������2�Ƕ!
��^x��%�?���~��_>�C�����׫������|��|&D��'�j*�e�Le��k��;~��@'�E�0��`�����\�^�1t�_Xaы�@��z�4�Q!��̀��0�ڐ�t:�Q��BE��F���2 �uG|���or%øV����A�5�@��h#LnV��.��1mX��\9K�.Ķ�c:�S?W��TF{
�E�e��O�l.f$�8l��|����"���(u�����l�?���D��Z�3!fݿ�ʘ����H  PR�Q�yώ�N݁7y�2�S��1�ۈ*�"׹��k*]���x�@y�������{��,���]�(r�w����06�>g���F�l�ߎPI����%��(�V�J����$0؜��N�47���Z<ƪ$�f]45d�G���f��sfQ����F�k5ǽ����)��-T��#�5*��7��d�wm�ƗQ׸s��Ŷ��J'�[�A��ɮ�[Wz�\��U���	�Y8f]��"fڲ�#���X���!�2rsZxE��Y�"��"��Iy�Ƃ0oh��Ȧ*柂m�����_K%ړ���!���H��3�}�j�u�o���ző��N�1k����>��Tk��/������M�!�`�ᡎ��!:H�����?.�����=�H��6a{�}� ��O+��̣<�� �#_ͦi�0!
�.<���x�Ʒ�)h/,p%�=��UȜ��]u�c�4����e�����Lu	�||�޿��OӀ���R����&�g�]��o�r4ix��ͥ�{/@Z�5��c����k���g�yz�,���4�plZ7�.aw�>�_ڢ�ɿF��Xmf���(��Y9���n/�l��5�%��ɿ�a�G���)��)�[{}M��M�Dwm7����[�l]LYg
|�{m�|�_7�����BEqv�-��-2���'{���2h�E6І��r��� N���Ǵ���/j�(~]faϭ�
��o<��.���Y���#�Z���͌,1ԑ�V���7�N
D5��F�z��$��L�d�����)��Έ���Ԑ`�lU�F��9���Gzt�\¶��Q�~�akf�U9��b)oKB��>�M��b��-�O{�V����P�%����L�C��c�d����iP:��iC�§��/v�>T���~lk_�����������B�y�衱�y��{e`��k.��=�#�����AN���|C�hL�����W��M�҂��IY��m����#���'OQ_���W���|��'���0��yHN}8I� _ ���J3���͸`�] �����������9��`K	���O��T����M3R���Rٲoǟ�sp+�?28d!$Ӓ�ٝ��(=v��\���~��%�36Ç��Gu�X}�3��7�B:�Z�`H��W�FPiq@�2)Vzi�����>�]v+��3��}oTˮT���4%F���ݧpdn��G���~��X��Q �bMw���
��TLT��}N+�}��VИ���IUv�\���}_F��0�z_W�D��������t�bQ�{	XE��@'-�o\�a�лGy�UJskP����=F�����+�y�#����L�'}�(꩹�Rv��|y���0�0'\.]I%[H\����sD�D_��X�ke��T�I܂�(0E�
,�K��|]fW�A�U)8]���4����^�oQ.)��_3$�E?�7yY !6 Q�  �2x���7\���t�J���hz�jB��\5� �hh�������F��]�2t<��bJ{ߊ��p���Btѹ>\�������̒�|�v�.^7���b0��	����#�s�V��37:/x��$�d�NH���T�@�^�"%U	��X�WK���XcF����$��wDF��#y����Қ�%�ز�I���1C��|hV�h�쫬-���>�tN.��	��G���z�D�ҫ����q�d�]��ޓ�k�[r��B{�t��P$R��W[:NT�d�	b�W�l�N��5���{�a�#�|Ek�D��_]U�n�7�::Nn*E�a��(Tw�9n�H�σ��˿]�1�K��,p�..�ݨ��_;a�`>�k����YS�Hmf�z��V`R��x�L�2�W8ǿ �{aȷP�
Tԙ4ϩ*ϸ����ҽ	LzF	�cs�=8>0����؟�N�Z�ȧ,�Z:�s6��̻Y���I�%�I(�9Q�Y�������[�8~p�Wܓ�Mh�s^�kX�QE��`��z~��w���]u-C|j4ȩ���*��qc��F Ή���p
�.���V��d� /{��Y�f��e�傜����YY9�b&p�-X����fg9��ղ|�S��Q���G���?8������j��~G�b��lw]h�a��A�ä[�׮��z�c�Q���κ�Q�hC�ʗ$,=�sA�+�f�������Ok1I '�݋}�����a�f�B��U�j�6B�����A�X��-OMY4�:��3������;�yٍv�<��KPh��)�
@��(��q_숄��k���mX��ސ��I>]�o4k��4iWK��!j1��U�X;�gL���j���&S'�Ȩ�����-��ʃ���$�����h���3��$�0��e~��
���m�Lt{��;�]�g���4�>���y\Ǟ(�jAb(S쳂�&C�)?[aP'�M2�y�iwV	�5灴��Z\qvG��q��������`o�p�fP��aft�E��s)Ί;bF>c}'�mX��!�Ht3?5��.�x��B����\B�*|Ԕ?zj,e�KH�\�c �
p�GV�{$����c����;����������BuXJU��pi(������b���=I��D�#�{V9�� (f	b�u�s~�O{��/�Ma([�}W��6�g��$w���^����Р5�j�uޥ�Ī݇���sZjIg_�Ѐ��~ebH�<ƛ?��U�]˃{���,���a�/l>�����H��څ����ޚG6��p��#�M>Q���Gv���!5�@�!�Z�m�7ߋ��Y�r��&������z�s.�q;����!�h?O�F����IQ�*��s�h�B�Zm��9��H��4�!��	�L&[}��0y7��}R���ܵT���9�;�Z�K��9O�t�M��{�쳥�(5y��{�@y;��@�f�h�ĩK��`�5W��'䄼�+�G�]����`?%h7x� dN�]ZfKv�Nc��7ukx��m��uU��^X�Uǁ��ȇ*���94A?j���+�+?;m��-<��}v��":�sB~����3`C��"^b&�	6_�\޴�PGzO�@,\wJ�:�,3PN�zZ�DdU-��q�%&�߾:�% �m��|0���QD�ۯ{e>��:��A�/�*�DÊq	k��
w�U�ǝ~����u '��}l?��F�y�Qh���w��(�9�E/&�*:��e���`R������FfB��黙�F�,7�`i�wJ��CC���t57�ӽӼt�\�Up���C[D�J+-$�oA��Z�B��������2�SO5��Rd�Gi�B�y5d��AB��|�5���/������c_�v��z-�y���o����}5�-!�s��������� �ޣ�P��a�+�����ot��k�>ʽ�h��Y�} �WO�*�C}ǖ�rG��_J�Q��6���n6��dH���2���Y���+r�X�+leCW-!VF���F���X�+��]��a �$�D����q����v��*2�Y���M���ҌM5G�����Ի���N�P2�1fIe���q�G,�D���|�ĥ��Gr��k��'�}Qꩀ��m�:�5]]t?Q,�a�4_gCx���wp�mB�5��~\�V*;f;q����PkB����͠��~�^�P9?�2=��+�~�A��tŚ���T�*��x�AI���;����~3�#��*�lҤ6�2����ir�,b�l��aT]A̡��6/�#,/�;���afiV��ˏ�h[��	��_�����uξ'v��<"���&EF`��h�t�X��ȟ4y���գFc����������u\�>r��q���|d6�	�n�Y��L���K+�G-�huU�+���L�䚂F�=`@1y)��}�Ku�N�
�<�$��5��?��q�*A���]	�^w��� )O�(�yVfk6��������;��D^?JCp*ߛg�"�c����*h
�.\EMb�>���."�
�}�v�����ǅ|1�LDf���%�`���~��g����!���O����]#�|���������R�G��,L� ��dCQ� ���-B�?�3�bJ;=E��rȷ5y<��R_��XI�{�ǳ�ɞ�EW-5l�����A?b��+��[:�j~ .s�P�o�v�a��m!�?�\�^/Ᲊ�Lyc��qGD�KЩ垫a{�Q�x�.�i�1����+���
���<��~���'�'��\N�Ʌ�]���u�����۽6}�3�=��U! ���﬜a���A�t5��{�m��l;y)u3S�RL �lYl�R�F���*=E���>��X�*���^��K�q�b��#(0:'�He��7�J2��eUWaom�FH�m�nܲ$o'��{�1HS�D\�h����3�!Ĺ� �Ѕ��٫P�!� l�ʢc�������g�0�Pz���5dm>���NF�j�!4W��Y�g��3[AP��G���P���a���_���}c��4Q	q.Kjd�C����G0�*�ֆ5�|$:�[��k�t��*<?b�>�֋3����"u�Y:V��!0����=��1���~8��Yf�� HC�����]�BT,��yG�p���"��x���7�W�(#t���݁#P�����(Ё��
��7��y�i���W��A��029��"�N]��L�d���e,�e��T�����~�;���������b(ޓ�
�f�Y�F�0��n�I��xEA��?|�Ȥ�E��>5(�k���[xiDJ֛�y��r^�J��f�˚�ԑ`����/���&1cv���=	��T����~Mr�_�"��7U����Ǎ�[S���kå4f,BZ�s⇛j���?�Lص��ۦ����>�v��f�bI��f�o����<!��F�i�zL���3�c"b�LH/a������u��Ь�n^�+z�Q	��w�	�X����u�5����,�O�#���knU}��sR���� ���h�T�&ybm/BMJ�r-�V���'#H���9*�X~�(�|Zjp�6na���� Q�n�)��"�j9%���~k+y>W�H
���)�5,We���'�eq�9�����8EV���c�\32
6*�FҞ;��C���;�L�����R�w_%�%�qy}�v��?�)4��(�"�WB�
�S=���;B*�fe��Ǣ��q�F �����y�f�4���x���$�M�o��.�@R��#���IRV��3պj��0�7YC���p���`�/=��	�#���PFy��_7،�N4zg�X�2���}j����nm�'��d�-���g� ��z�y�$�m^h�Ӯg�&�8�zW-�sy�D�[���ﰯ�ӍlѲY��k�?z�MC���͈䛐�d��gs^���URG���S̢�*������U��q~���-�=�<��\�"�@�rnl���:�q�� �T��N@Y�ƣ��5V<��O�&ł�yJ�6��f��Y(�2ǳl�F03k��2���.�5F��<��Ai��J��;��ÅRQ�3e�t��<j�F	�%�
ɢN�Eʬ�S��ٛ�wD:�]c�n��R��K\#�a�AA�
�g�;�n�|lG7���|N�˩ 9���!}�Z�@�?�,k[��i���	�� N��`}��5Oh��Z5�r�"�+L��|t���A\٩�#��=b�y�@Za�"�JG�Q��J�O��g#�z64�`b�מ+e��Rp$ɸVձ�_��1��E��
���T�jKf�Rz�Gݙޫ��
�!g��^�� :d��8�S�0J���ѻ�eԕ���;x~�Lb�%��Zv�Ղ2�!޶�r߾��R�y����0����S������s�*��Nt��Fô ��0����I�d
!�Af���J�p����w�}De��u� �>�B��n���C���rj��0P����u���~	�V�i�� wvT���'��D8�a�i[��Z��2�f��د�,�]��J��h}����i�=���k�4�u��^zIJc	-�ۧ?���Je��� ��?��u,6��/���p��k�䨨��9��_�0lR�T."���wy)T D����ًxC�#����^c6�F��5�wh80ŋ�(gm�&�6ܡ֌�F��O��i�+�Fu�|��c_Y�.�?j���W e_G���U��%��0U�������'�=��Q!��:��0к/p����h`�<)H�t�Ó��o���8^�=�ZԚ�6�w>j"���;`��%'�MjBSP;����G]Ea't��"X�U@a���Ӫ�C"�RrD�q��U@�:���~j_2/ $ ƥ��c4ߗ�yo����y
f�R~O:_�]�5TK��<˰4i�c���&,)n�f����m��~�ߜq�us:�z\�Q�Z)��t߻s
��`����fڂ� ��4|�8�㑵;�T%P�G§=d�00�����i��[���=��u͋��Au��� ��½�^Y{[��Ǧ�}�K���]�����6&�m��jI(U ��#~"�O�h��o���?E�o(ik���e]f8�*"'�2���q͸���m@�L�8q��`�#��XB����'R�K��h����q��Gػ^���	r�tU��[t���В=y��'G���y� �����u�R:9��u__-�r14_@�w�0;�v,{�� ��W�'�����g�r�7�T���,�-ͷ�YZ���k���m���ө>7jB����5[9]C���I~���ݡ��#�{��n�e��w���8��I_���c9�^ze��"3b�Fo��X���Ы�Ko�[�>��l���Ag��z�}揺�o	����̓z���J�<L0�agC�h����1{�AN��A�~��g�y��E���e�C޿�� >�Hn3�WE^��d����i6ŗ�<��/��Bе�А��4�̤��]m�M���X�. +t`��y�Qa՛ԏ�~� Fn?<i�2��#���������\{$�lc �Yd�Ճ^`@aq�����p�.k5��?]���ޯ9�Zq4'"�KC,���L����Hw+�Qz걐�L!��OŰ�V�Pnv�sO���ZS�T*9�^s�Ї�Z�K5l\�~\C�� �4|�������(:�p�o����po .z����	B3��6G*w����oʬ��)=��r�Q�~�� BG$:J�a������п�t��l����˵�[����Ea���Y��-
��+1�r;��m�@N�8Si�_c�Aƃ�Q�(CMq�4":��z�#��2��ǩ�����#�0Z�eK�M�.�09$i���|6�ǯ*veVա��O�$r2��r�G2O���t�?T����k�lcbD�. y{	`�p���w���ۿ �,_�L�7���x&�v�e�ʷ���z���L�~��Tg}�pp�c+�P�D<Ŗ*�!�O��$�fg=Ůq� �$d�-�L�UP�ap3l�1y0��R��pBduv$)���5�C��i�/L�`��)UَZ#��_����j3ñ�",��|�W���`t0��]u���)�g��N `�\|T-G
���P�����cu�cjl��|���m��&һ}�0/R���:�M�|�\�]�����z��%@xw��f�i��t�aq����=}Q7p?������_����y ��jȯ���l��v5���5��sKbb!���a&���L��0���-�u�BX�I0��G�"�/	0G��H�(~��z�/��^׈��H|�`�2&��-D��<���c���KHBE�>�i|�r磛k�D�����,~s�
JOBE�`�lա��ѩj���*�r�?������;���3yc	2e9��A�lLZ��1���L$��")�Bc�o69��~v���hU��yYm����� ���pEg�Oa{Db��	D]+�&a�"�p�Cα����GJ�߁��.T��<����Ț�n��SͱO�V#�(q_�{�u'b��߲��AN�p׿'�:D%��G�f ? nM��R{sd�&�J�s@I��5���k��`�q�L|�pn�Pk�Q%�eY>��0L	��X�~��:���{�E�B�K�lt���s{|�r��<C�j��� $�)ʁ):�U�~{+!zb�`�r���@���{��A���+�V*�@��ܟ����>�}qZ��F�R�|
�f��j����a��{�Re��5�6�LE����|�E�a�Ǌ�w����'}��D��~Z��4�=n�x��.�о��{ˀ	�}�ђ<�<��m��\��l���S�	L c�*[�������: t�7K)g�H���F��Q��A��h��Did���Ah� ��@g�F�DѸ�5uJ�N/9Ы��Y����FO�#7�#���<5�����wf�O0�9�2������}��iԂ�f�r��2-��j�ɣv�}�x��;�"l�R3���V�r����/��6"@����G˯n��%+�j�&�x��W�-u1��x[�]Wyx��@�Ia�iP�Y���>����������j⟬*ƚ�9�s{���D�g�u^hĴAUh��t��dj��&�����`��;��t]it�������FP�pfmy�~Њ� ���J|	e<X<;��F����֕@Y�y�F��r���hϲK܍�A�݁�N�\g�H���S[�2�� ���&��@����e`�������� oy��AC������"B��*�_+>Jq��_=��u��l��sGBZwT��%8k�X/��RSznа�������0�KAT�S&�xtw4�A���;��������}����1��o��Ε:���S��i�����a�c	����0�8�9(���R`�,��z5H��W���պ�p]������5�Q�߲A �K�F�[��t�Z��%T���JU��~'�n��Nz���h�@Q*<;A���B�U��
�ː��e��{!�*����N`�U^Z-xܡ9\�jr|D�2	��$[���@��{p�KC����2z3��ظ��<=�*�u��a���X^�OE�����ᣅ�ː�ǟ�~�H覙��s�2�-)���YN�������9�o��B�!M��{��W���{�5�9����Q�/��M=���N�o!fJ�#r��Q�IAAD&i��R��Qi_ ���<��)g���r���㹱�.A��3��k�� ��kW���6v�-] ؚ<���}�W^hI�+֧����]�d�����
n��G'1HQ�i�*0Ob�I�ӡ���@7���{�%�O�\@1��2=fF8�&��d����}�E왜�jL������#~�oߟBd�w��G^MB�n�(��5�J1���HL-���EqA�B��I^���K�{�$ʤ�(Y�ğ���n�e���8ㆬ
�Q"Y��������^ڃڊV��Z�����^(���i����Z���=ג��2�����
�#��H\���_��d�T40�C�	��V�%!8gD���5~koY����$��ˀ�e��e�y-��Eh��y(��!ɮ�a}5{6'5*n8�M\���Sޛ���I@��;�NZi3	��[���:�Rשչ+��t]R~y�L�3X�͉���0?I��X���;��%L6�zo��F����y<r����2��3�|������j�*w����c��B6����$�4�eu��Ũ��!A�x��9'��GUN��m��_XK�-ޜ62IЋY�-s-�{{�.Q�H��:�0	���O�\_��M�l'?�V1pe��;G.U����l����v J���R_���!��k��Y�ި޶pQ詩:߷��1/��	t�4�Iw��:f���{�^��m3��hS_���-���*���Hp03�X͓�:�C�w��;���N�x�B���xa�������vVӪ�����_r�\Tg��Դ�,f���V��/�۵�M�n�x79g"xpk���[DB�Ϯ[�������:��~wD|���ծ�ׂKg��)E�=�_7����sԳ�H�����8�o�@Ѫ|vb�S�Y�i����,����<�ÇǢ���Y�'�.q�ah�9Y^E�!���>���{5vغ�]���ͬ�}�k�=/M��Ň�g��x,7,&k���&̮(��zk�R��n���sU��ͳe.o���<���	�~��⪗�i����,f�����v�L�	��#���<+���H���\sf���X4��KG��	C
�/U��o9�г��e;�%�����1AucC��3���/z�)4%�-a�M)˔?�� Rm����血q��fy��[��J���۟f�P��Z`mZ�8Y.t��vc_��Ib_�R]gɭ-yC]ͽ�Gڊ�����s*�_��KXaM���k�L�ه��6Q��ܬ���NRae�C�Pu?�8�#o��d��ϼ�ڂ��˭�Ƽ�Vd0��w�|�P�d��Z�L`�U^�r�i�X��	�S��~ARy��I�ƍ���J�ک>�s�H!h��kƹ��{UIj_��>T�g@z�Q��G�rN�Io[���r}#����z�����J�^uO�'�*G��GW�f�{Ͳu�U�����b�����e�GQ2�=��.>��:J� �x�H�����wF>!�Yv%�Yp�uH8����/��=��9��K��-U�ٿ}�w´�vbX� �O�����q.�o�v��W�o_��mN�Ζ�t�ԄT !űܓJg�W�+���F)u0��S���L��\���{�H�����=�oMc'��4�N�����	!C;B�t��R��t�HncM���,�����7as�b_�J���l�J�����	@����.�	�3��d#��C��[ZOD��6�$�f� qЋ%7T�r�D�[~7�����^฀�L�Jy���b6V�5��`�w�w����Z�I,��⣀X�G2O	"�J��L�J�t�8J� "!��������������:��`U�Y�D7J�����ݿ5��KUWI�̱Q���sU_�1P��0wK�!���=���e��C��m>u�D�J�����^�Ϣ�|a-�������ؤ�U��ٳ��"��[c�8�r�C�]U�
�z̬>a��o����Ć�cy�g?�kr�r��'��~��p� ��b�����-���8Y��;������-l�L�wS/q�>}^� v���� \1@�czο'%�ױ�����P�-{���qA9HާR�DN�g���OY�1u��o�9?&�a���П<j�@�rk_KWYj~/��_��;t��*�)��7�'"'������6�ߚ�5�v��Pzk���L�ɭQ�B�4�.6L�w�4?��~~������Z����g��+h�5I�=jn���(�֎�����6���'�O�>�T��3y)[m	K��;ԕe��f�&����Cs��b'k�^8����N��S(�,t���p*�c�w�n�)� ��I*�kO�����'1?2_��p���c@=���~����P���h]�z��7k̕��,��AP`y�S��z�\�u@T�n�/!
�&�ylXW�4�
](O��k+���G=/hv�BBkX,
MJ�Y�^��%��9���6�|�fN+���u�� ��|f�U]���o'F���B[��Sz�Ϭ���z��N�����s7H<Y�s����@>��B�/Q�:M8l ������7Z/��F,�����V��#�3�%���3��h ���^Dܤ����Z�~��I�hP2$WV�����Љ$�~�֡��ّ��cl�ky��@}|�V�=�/�U2u]���>�"(S��56�ڧ�͗ҶU��S_�a�SR�|4_���D��Wm@g��Q���AD)����!Dk�k1�����gD>��ń jWN�����iG���8+q� �De�*���y�� #�!H��+����-KjV�d���r*�X1������Ԣ$V��L�|��qNeV9���2|�z|���HU�-�<䀛�g%�zQ}����dTd��;.+e2��Ig���;�Q��l�)L[4��ۑ��*��~�A �<5��*�0m���-�N����%�ԣ�|�s����w�^Yn�\x���;� ��,��'����n�G�x�aƧ�g�r*��A�1��;�Eԏt�������)�"N���%\�B<}�\oyo^~��ڸPg&ǋ*�jb|�N���R�����A� TZ��a⊭���ۮ[;���D�U�S�-��+��uET(~v��t��-�x�l��kؽ����&��N���<@J�4Y ��?�	Z#u~U�O��k2�)����7<S���k׈�KIquȧ>�if�{�b�%A�N<%=�ґբ��<]���} G��E3�P�Ͼ,x����:]�W���?��h*�w���K�Ebm��arx�>}A݇��u|��A��4�ؾ�Fr���{c���cv�(<���K;O�_vy[�g�F*S�:��nJ8��
W;qN����5m��������j���@+�.[o����z�)���p�G�2���3L��]]B���;^�������P�q���"$�w�"co��0�~P���! 잳�l���7�>���%�pu��}���׹88x&��t��P�� P��q���,�����^���	J��A�i�נ���s�i����E�j�55���[D�^!��MA�sȻ��Aد�ә��;���f��1���_*r#�s�Ҍ��l��i�@�*r��{ԴM�	\�3��dOผ�� �v�i�GV�Z46D�:n�ZLs��Q1H���V��c��y�a%����/��᠑Չ�Ԛ���b����W�(?�z��R�e$�^Ǻ�@ft��Es:�B�!h�!&�{:��Y�V��n���a��!�;t}����5�������Rj���� 8��
��i����M�����S�U����@@���[w�uj��&W��u���E{��~p�n�`�������:��ײiϪ�� r
eIEb���y��: r��{�E���82sE0��8&@�J��(H�aT@��@���q�$ �b���t�A����6�dhr��9U����_��/��Z�.ƪ:g�����g�*��16��#�>B�ƭ4O](�D��y*�W�s�Q��Es鄉�:W�?Ij�W����������l|��#OU䢸���� 5N�Ӥ��Mx�!M n
����/&&>U�F?�Y�8�>�	��5>�Hf��v-t���Cv��u�Dɳ���>z���'z������L�Q
�D.��j������M��hc�����%PN�1��I>���^�׊q+O����!��|��Z��dX4����� �Z����(�N��ڬQ�����vv�	�j�A�ϡ�fU���eUA�~''oA�.�$u�fs�ʇ�R^/-F>�����Z���A_Y8C{F��~0���.�^X���@R�Hq��H�C��&��7�[����(˗�i��� �j�?P)��ZCQƞ��4�F"�͌��)��1�_R�ߢ9/��ާj��C���e�Å8&�������G95@� B�I�8��4Lw��|� ߆�K{}!��c/���A��-���N˧�xl�|>e���U�둺@���	����.\8���֧�t�g��`��kLl|��8���A�����&�Z�m��q�#7��E�86�н�����PY����>:o� V|�&��1�c[�����|�mBڗX��:m}yױ��HȒ=� Ś�q�}Q��uh�x�xg5tv�Ә�9/���ve��VQ$&n���8�X�n�?���qA�6�+(7��6���2�Kq\:L��1�����tn��.�$G�����{��)�/���F�MT�-�����E�s���pB�^y�,}
�g�o�̺,|������X�N�;����]�ƛ�HJ�7�ThtMAr�n/���j~�~4����P(����(�t�p%r�vH�@>��~���j���Z�=���:�͔�A�r8�H�@�M�����9t��������?A:o��)��ǫ����zty�u"ȴ����)k)c�S=�HsG����U�Li�N�����Ȭ�e�B�dz��5���ª�w��ɚv7P*��G'-�*�� ٧����n��c��oe������4��+��<���s��*�lu�	M.u7K
�zϹ��k�d��x+I�.���bD ����&�Џs�0e�u��N���}�KA$s�x�	s �v�k�(��d4�&sG��u6/>q?n���:��v�>0��� �����Xؗ�M��~̧�k�ae�b# ��_�����P^2�R�h"��l���S�ڦ+�=�O��}m���?N� �-�vay�*�����-yF���!|��#Ӑ�_�����<NG}���AX����9����C�&A� �Wޟ�(��:7ydw`�Q���RՕ�gzz�\}�|iq� �����$��@z��\�r�U�#ਝ�o�������vY�G�~R���@i��;s�별��8��Ey�]����/V�|o��]�$�����+®~㠲6�j�w)����{ޔ(#�0��s����d�����j��|��N�/�nϋ�W��ԓ&��j��WN�� �Y��Křƛ ���jεq����	�╫�"h���%,(=�0iw�Ջ�H�w��#�������p�����g���C�U�]�ۖ��{�QU�j}=�r D����Y6�9է�Sչ��%_J��̏ �	�%�,x(����[H:ICtS�&��.�y�[��s��_�207��W��S��f�Hbu�.�OD��Cn�#�* �����^���R��Rl^�U��$�P�{.i���W�#
R����1UP*�<K�{46Jy-{�����"�����zQ�~k^��O�Q"MZ؁� 5������;���:*(/��C��k��(Q�g����MoJ}gG���S�}%L����& h��AR_���6�__�vr�RP*,n;�s�O��MM��9s�> �ȇ��������W}d,"�#��Tlr��]�ڰȿ �ʾ�N��.�e��N�$�?B�?zT%[P���T{��K,�7;~K���q��-�������������'���ؓ�ҷl�������h������cN;NןY���iX,��o���^�s�JYӣ���f��n$q�Qy_%�ڽ�t(jjEU�%o��u�m8��\]�4�ƍIe�76_�n��6Vx��Im��9|�[�b��3�S�[��W�,��p����A$Ҥy�Ło���K��`�X _L�rX���t�h1�����7�8Y]���&�~>�섋'B�]�k�Ȥ�Ak�M��i*H(B��*�1�e�!I��7���bV?�Oۓ6�^h�uF{Bq����	�U�N E����N��)p�6]�����n>�E'�8��S���!���>���۞[��I��EWE�"��Yx��Nۮ�>d�9FuG�ĵ��"���yu��K<4<��%���g�K����V�Y��S��J?��lEsI��v���'uS���Y���Vm�G򷄽�sm>[@9���ѓ�9|���GWzT��)�85S�͈l���D�����:��,�r��'��%hv~�n�Y��4l���Nhp���\�l�Y�� �'� _8�#'�Z�/�#���ا��9��[�p�E��v/FG�7��>fe˕\OJ���ߟG�xNMJ��e%1ڃ`'R&.�S�`�B��.�Q������-?���i�w�oD���?@
�0�x>ٙ5ݏ4�(o�m�{MB<�:�v�{�κ	��V��Y)��k<����n��o�^�K�B$���&QFs�u7��i.����ȁ��吢�6�!��$6j�i��،QX�X<:�� ����y��l�~��gAα��!�-��_����z+l��m �B�?B�*��Mg�n�:ru�˄��n��]�>^	N�>�f�����+��uҙ8_�''�zW����&�]l���nu��Ǔp����;�ޭ�F�|ҝ�wϪ��/�m���C��L���7���Y)s���'�YI�E���0������l|�!2��:���?{��q��sk�r($�ԇ��48�~uJѕ��#�p~��T�C��l��;͢���z!6^G��9��҇�:���u^H'I�H滤�J��s����$7.x�:?���kI���y%�9Зڱ6zQhf7�.���L��F/���/`FjQo����&�Dy[�f�_I�O�)�]ob��߀����F�6N���]o+7{�������,���g32���e���/f2�"$12���yO���=	�p���U�Z�riv8=���2i�2-��[$~�߱���]��p��BFQ��rH� S̦ӓ���	GA��壟�k���d��- rg�p`WZ�DMsE�#�*����f�e�ꕽ
ܥWƱd�T���)1�(����7T$L�����Nn���|d_��z��z�����v���q�1��NQz��B���k�B��]���G6�8��C�J�A�{I�y=`k�S�A��B� ��w�]�?��/��0Eo��>��e��0��c���Ŕ: �;+��$��o������O4E�먼=O�6mH��<��%������%+���0@_M�	'��M�;��?�I��p�$ǧ6�F�	� i�]Œ��UQj8G��с��y@�#֖V�����z4�P�y
t�g@���q���!�+�S�N��y���SB�̂i����]��2�W&��خ��u{%o��x����;E��ԣ���R�O���J|[�@��P���Y�q�Z��-��d�C�ss�u�-�Ps�L��.A�Z8\��g��Kb-�^fj3�,�31��L3��bq�z5�_q>�t'��3 ������,X�@&[�Y}�^�Z���.�7*ڡ�aa٘?��&��UVeFa�T�.Hfm5W2oI�����3'#�_��LB�\�d��rҭy�6�4��{pN��C���{d�_�G`H�X~m_&A���2Ǖ�fq�3)���,�/��.�u��	����.]��ܩ��+�u��՟Q�˷T|Q*��`��(�&�������(����`���9��{�F����Z��X��<�����=���R �u������y�*��:$)	�o�Q�R	�U�����he*\����>�Q���c;E(ݥ$�4)�q�{L!gŁ�͛	�E�w��D83x����h,,��/i:�A�@�w"�]�u]�ׅ���63����|ݾG�,������欌����B�A�]���i奡��^�A_������3���ѫe�7��<(@����	�9�Q@�M"F��܀[*=F]J՟���I��׮a�1N�%-:��T�䖿p@�#6�v�~z��0P���߯��G��f��~�"e0�qFSO�0�Pl��ˤ�Ԫ��`$�� �J��S?􍣀�$W��W���T:?O�É[Օ��D���m�!}�-��ֿ�[��B��2#�9��>�g� �n.p�(g��<�'����B���0o�%K[��a^��2�Sv[���a���[ ���Y��ֳҗ���MuB{�Sq.y�Z�' ������:���Z��J<§+O�AUZ����Q8i͌����'p�wO�_���~,3�N����@��a��%$��/�vP��[��u+O��i
=��r��ڧ���D�r�mA��#�-�B���d-���*��S� ������,�2���L�7�%�����S̩���C�N Q{!�̯���T�e��7�~�N��p]�ج%E��I�pڀ�jG2�����*$��]I ��$��E v1u�<®��;�\_�E2lC
��vg��\C��K�;o#pY��g����g�k�J��9X�j3��� E�\w���g�*�z]8$��"�bg ��o$)�Lʐ���}�AI<�i
w�$>Y�ʰ��}� ��:��?:|�=�ϝIN�ݏ�D��v]k&A�d8E>�����|I�͋��K<h�v.:�muf%�:�58�ȧY��b�6Ԁ+<du[�x�q2��!��[W��iB�<�� �iݮg�����ӂm��� wn���ɬ%�\D9��-_]O���h�uM�b��� /��Q���_F�$�!.�jZm���w����_qu�K�ɡI
����	�=��,��Q�v���p!��,����"NN�~ѵ<d� ��RAx���=�����k]�ɇ��tt�
+�뷸�;�S=8�L��@n����T���֋��R9�u�#(��M��j���T#� 	^�Oߡ݊�C�=�i#�����#Pa� G,!��}��7��~*���������>�-�b ��:���.j��FeoWQ�j�-��e�"[n�-���Rn:0�Ӎ�^�$B��^�(���6$ܧ�V� ���q�t��b�U�����pokK9@�:*�j�������Vh5���Ay��)��n3�X��^�iZ
7p�J�ƚ\P�A��jƢ�oc��c(���6��9���ihX�V9�|c> �M�z��3e����+��8��Bn#�w&p�����Z�d�yU��,������a�'m&���~4x�RO--�+�N�3�N����E�D�"��j+�D����j\�Bg0l�=5�(g4�ts��+�>��2�Ek[�	�v�ӕ�od�*�L/��i��&�/�f��;�p��$�f���j%�9��
"`�2�duzm�()m%q�4�irr��0lX��{8&��৵@�������ڳn�l�2�����+WϾ��d}S��[BK?��o����Jl��$f)J����嵻{��C1�K+�*3�cZBJ����@�ì�<���89��]C�&]w�4��Z͌��\���cR����E�~f�0���U
�������BPS(�cRj����-/�dBAQ[~���A.���4��*0� b���w��0��n)�_��K��nvjN��%�҆k�>
~��>7k�S����~q=��V4�Ք�;<�����ͼ�f��#��t�#�eU�����g<�T��B3��Lj����aM�' ��6��k����/��o������ �Uc����r>	��P,~�罤�$����G�m�r��
d�$�/I�>�=�����B6�0R)~�����(�ˋ�l�S🖟kY0**hU�
X�%��e�R�(�K�j�>�,ml�P(����8p���4$r���mEd���x캤�Jc�1M?{.�VS�8�(��+ �Ճ�����6Ȋ��K�.G��}��\�|������uP�(Gw����?�v��l�X�ȧPTV���sf�	7Ɉ#z�nŗ���C��n&��ОH$w�]~���P�Dyt�w�C����g�3��t��>f$T3k�9�A��9�<8!R�R�gpf��:��Lu��F��:D���+�����u�����W�&�1&���6C�)6���c�DT	w�By��8�����~Z�z�!&��%#�]���$P��w���ؿ�I��/�� ř9�A���֬��%�Z�{PJ�RJ*�m���*e;*5� 
��U|��P���\�&o$���<��a't'��.׿�����vγ|�p��ˏ][��>n���FҒ�2�z8���_s&6Qޖ���w�we�5���u�"�v4��Ш�Q	��T�v�����p�'�]5i
���q,;S��e����dD��Zy/�6%2!���˼�|o ��:y~$UG�Lo�7�[w(A�	[��ʙ�	�A�dX	�7o�dOqԨa�+����#_��d0��[]�KNÎ	�&�8�39���}�gl2��|���|GM��Ʒ�*�=b���˾���^�%��޺lo{#/�-�$O�2��Q��݆ks<
*D�^�~�O��T&��8ny��c=t���Lv��QH�^�U�f����w%<���<��δZ���<o��w�.��!)ÉR2��B\���݇�SsAƾmf�Hې��~��Oq` �ѯ�ߟ�;�x�!]x�	79\�������d�Ƶ[�Hg���s\��:M��D��g�R�<y#�㰠(|I�e�,m���b]�T�	ŵ��2��.�}�QA2;<�n���_�Ar@u�9��Eƪ-��7��7��Ѱ����%ʿ�i��DK�l*MH�i���"�k�9V~�
;�3B�o���ʖ~��L0��$��L�]sȊqa�/?@&�؜�ޚ�9< �N���GM�7�n��b�$Z�� �4�Sϟ�愘(��*X��aO��?r�PK�EFTJ��������!��O `��
O�qUd�ۍ�W�5�9]�b�LR��G�	ܛ��Q���!h��o,�|-ކ?��@|���5��[E���a�v1���Q��*ʅ�-rی�KC=���@���F,mzE٨xA��ī|���p*�F��6P}㇗�P�_\1���������N$�k�B'���a"w!+�k7o�8T�P���V~7�:�i�U������ЉUO�p�8������t`�o�Í/I�+p[z�C���7���'@��`���cΗ���3Q���D�(�*1ݺ7?"��[���O��p7��U��H��#/Hp ����3�q�<D�|B������w䳦F|U=Yg����̚�\iN)-�b߳dt�4?",~�	x�f��g^t\z<���-��~
�]��vF1�&�B^�|�_����"}��(Jf�qqwo�6��j�,�qH����'��I�.~�-�= �~����Ȧ��D�W�#.0�w;���Ӌ�07q����������)w6�־��($�M�������Y!̰3]H`��R��0�;!՘�N� -��;�LC�i��g��_�Na�2=rF����m���-<�&5�2*D���������;o?L7S�F����p�F~�0Ʌ������h���&��#�!�թ�M�_�o�����1
t�9�,��=R����_�+àl�]P����{שZ��H(e�ȘC�x$�������M�����<� �^��J��_6_j���.b�Q#���۴�y !E<��<Cf���#��{�<�E�p�����ʰf< ͊�˜/�S��HNS�1*�P����R���������d;7D�~�Hƒ�9) �w@��[8��ҧ����r��Mya�nٔ��i]�Br,�'8�<�y�ϓ�֔�;����j���V���`?#9C�ÓmV?�@QA4J�n��	n��Gc�.aw��,D�إn���n���Ƀ�=IW�P
��?�b�$�l`�W�D(g�����E{�p����s�Cۆ�|n��,���e��tDqq G���[��=�0S�뛋b
�y���m(w��R��iE]��|9�i�9�j�:Y��3��Q,If]�t�%�q��T��Ɂ�46�w{��mvK��0��5�0e��:��(�c�f�����Q�$�.�2��E�#�rm&� )+�\]���߿ϴ�W�A�`����*�����^���2ZO3�>h�U��K�������K΢
�T6A#��8�.>�S>�9�ӧ����B	SW���aH*�V@��N�t���X��&�����Cn���{j�C� ����zv����)_m�����n7X�k�3᝻�����L�y�8*8j�x�DW���E�����y�na5*���2�y2�ij���_�f���c�qt���I��6���f���S �Ct���H	f��m��δ��7`%#�e��־��Y���5J奾���)���}�c~�!`�	5N�������EƢ��?��d-�c��OTHUeW��G`���Y�� ���Rq2��<��\���
K��!�֎��i_L�Fk����Rb�|f0�?G$�����ל����E%��@M�$7֕(g 翲��^�G�d�~��BsBWT�H*XB��ڭ̕h��f�5z5% 
� ���7(��zRr� ͅ�v^5A�]=`��� !�grA<�!�'����im d ���@v/�ε!�kg��ȡ�������3H8d��O��ѵ�(	��4�D�s.b�M��
�D�l���,��C�zγ	�����郞'+�	�fL�}s���*�����}p��?,�&����T�w��f1�N n9�:8�N�?w	0�\��W�
P���Eg��@ß��m����Ⅸ9�~,|�+*I�T0Cҁ�<@�Z�����G��a?��fDٯ���ֺ�=��2$�"�$�L�h3Y&��O1j)�{���ֿ/{�!G����1���m2�.�����o�#԰]$ې��/�C��F��{r݌	T�͉W!ַ�'��)��A�1��5l���x�U�L���fp��-/��4�@m��6���܃�2�����'|�x��nm�6�~
S�轗�s�K�@6�lLu�ԏ#�9�  b�yzm	Pa��b�� h��'w�Hf-+I��j>�7�6��R0�T���œE��-BD-9ņ�5*�`-dVW���P3[+}�F-#1�M
@/=є� 6�B�_z\�{'��`�������j�:#`X�d`�%*E�	^�z�)JZ8�
 ��C|�w��fd�G3��R-�� ٽLȗ�	ڇ�����N�:���*d�h�^דe�"_���icV���`�ȔKX����"����(�h�Q�"��xBsY�\��P�~dw�^e��|�SE����,S�n^:����3mm��$+���vzX�E���F�Ov X8�ι ���45��O�e��õ�d3�G(�C�I�:c��m֮!�P��\��5j��M����}��o�=��
d=�9FC���"�]��)�#`B���O���,�8�z�;���;�ȁl�q��D�̲|����[�A ��������:>�������c��JK+Z���� 0�-���Y���Ϭ,� ����,�}�\����}� )֞�}�����������
P.Cy�W�K��k��,��v;Dz��M5��w����E,�"����f�S�|�" ��?���j���w  ,Ew�pml�`~C�]���Ba�L���z˷�g��7R��o���k�t�e�e��ۃ�'�1�o3A�� �H֝�����"��7,��n�[Ѵ=�I�E͙
�"�{U��k��]sr�qS^`�~�r:�>U~��o>iV�Di�+	���LO<���4loe��=�hL�9C���ٞ �\u���?����@��!(���DKuI!���򲪢���@V����Ϳ�௷�� ��w�&�G
GQ]�o��L�{��|�����^w�j�N��[W������bs�"��`^ 5���k�Ji�Z�h� F�?nY7�_�F����ЮV�@���-W@�;Fq��;ia��~j�ϯ4��v �f��jAR���/��a}A(�Q��&���!��|�u�M�
>6{��m5|�du�pd����
1��] ��A���鐏�7���n/lt���|}<�7��O�|�Ŵe(��\���@.�H�Ȕ�L�Yl#q(�.����m�@�Z�2�i�:2j�ζ�>�fBy>#�X����}fT�p��Iv!�Wˇ8�OUz� .��u���$�a��Iݗ�Y������~|� ��oi��fQɧz�Wm��X{U���?������XW-�����^ܳ>�b����=���y@�Mm�	j�i`{)�olEr1���&7/�6��*�2���+�w��}|�Z���@�w��I���F���[�ea%5����pdgi(硐�ζ�F^p�һ H����������O'< \�U�� 1��`�0���#�O���?��Nb�1=0��Uo�E���i#����b�"L*:}q�����`��6�г����8�{|�hw❴��1�8��\A�Z����#��K%MjFAq�L]&C{�}�$�F`8�埳��R�vf���Y��UJ��!s ���p�z��8�1(�E��D�,� </n86�t5�H�~�pfN�|�q/fk(kSdޅ��P�a%��?�e��qf��)D�.��<Q�X>h�X>&c=ٸ��X{:H8/����㏸HKב������������xwD�G �{ԗ3F��ڏ�o�3Kb��o��K�H
�Vב-��K�,����Pi�A&�b��÷��Ϗu<K_�K�q̺��S�l�޻�9OՈ���������4�u���颌��V�x�\`��Hz�wF��uO�������؟�[�d���i4�/>6�惘�Qr��pȪ��r�kౡ�(��kgb���}h'�ߊw��/�M5�h�ixAw]I�u9�Zҝm����D�%ŭo\)S����K���?�t��	����˭��-\Y��9�t���<㿲
+��+n�=o}������er�Y(�T��moV�)��ɠ>4z�]�Ԫ=�H�P1����y,>���n���(��+���x;�Bn5 �*rn�
Z��+u��_`d"�'�,s��C�(���5�~�ɣ����Nem�W�����5m<G���TI�x��=���	تwe�Vp�;S>�֢� +��n�Jp�a<��1�v���0���oN/x���@D;.��8Ca�|ES :eߑ�f�?���(�_zI�Ɇth$Å��t�k2*d�Ζ���'��]Vti��x�G��f��|(qu2�7!LN�cmlhq�,#H^�b�����B��C�48q;���^Fc[��
������ן���&{]5X�O��V9��ڏQ+^7{�J���=%
K�M�x�w۸�x�p��@�o.����4�b �DT�-�'Ʋ�M[�<�u<��dp�PEc�2�%����-�(��������s�{p�����[ ����yY�"�8ye�N����^_���ɻyfI|1 N���7��7��ί4/��0N��p�����~��{}���h�i���Ӱ�k�|L�d��;�F!P�uߋ�p-����zCgI��q[������`y��ȹ�+�3��3���t7���.{��6��
�w��xq��J`V�
h\O��t�ֹ�0��S��]�Xb|��Xߵ��ɼJ*���n7J��3���QI����ڱ���ޜ������?��W����^�yt�=���ª����ǲ�����<�M}!A���#Ul�+��^Ge3��{1�� ��0�g��_�8�0X��?��Զ�bm���	!J�9h]=�����k��&?��O�d, ���1� ���6��a6L���?�o=U��2nl2�pP��h�x2��Gb$|��/��D�y�I�!#"1,��7H���9�T��H�A�j �;ί�6��v�>M�������j����c�$����g��4����-��x/H��O����"Dʥ�t@��q0D��5��?}������c~����#_�)QG���9q�}�9��·���ќ��z��p�!F��j���i+�z8������S-�	t�{K�a�3�YG����x@��n�+�#���A��X �?C7�pZ��S$	pySC�|%�+�� ^��?��Z�8\?LAG�~�a�!���k��������y��x��+߀O(��s2�����u��o\h��0@�2b�ۙ\������x��9dq �"ұ�x<��5+�NV��	�v�9lNSX�� �@7ކ�S�>��4!���7; �Q��dV�F���y��c5��d�<
�o)�c�!5}ݡ��,��8ׄ�_J�$�5�y����\��)O0Q��↤b�~K�����N^pm���VT1B1��!�@�R�_��2B	�e}��T��1/����8Ǯ����r\��(+ �5((�I�4�n����i{R���Ձ�ޚ%� ���*���~t�	�t� �sdj@1�x�'#���R��c%�_���梻��̀v6��Dy\�����3mm��u�"y�m2��?)�f].y0�Q a�8�j���y��ZӠg�=<U�փ�jc$SS�=��A�ǁ���i<�i�W�2��] n��ټ�T�h'���mX.�(8���o,����3߾at���Sl� ���X/3Fݏ�V����«����Ҁ�H���[��>��3c�.�/���0y`���?�s�t5���X�.���500d�1���[7[��V[7,t�Ǚ$8��y�gs�hŕbƶ-tiw��sve,C�^���!��7�����PX���)��9TƕE[AS�X������~	��3��;U�%@*f7�?�\(�����^gCۚ�$ ����d_Q0�'��>Q�ɯ��dC�����kD��?�vz��g��\��Ji�+:�z��x%�T��_ +�&�@9��2۰��r�#��_K�8�P��7��.�0m�w���_��/���'�e�Y�d{�䍜$gDQ{]n��m�
�s-@,gvt�\el�B��X�c�N�ݥ<͏����]��G��������L ��|�����$b�Tݝ�c�3��6~�dK�&�u�������ף�(Y_���o5_���7L���]�Y�1\��^�Ȟ�	ѩ,��?G:'��>��Ͻ?�d��M��(>o�F����YM���@"�'��T��]�e�Xμ<���R�� .m����X43.��im�!/�WGǙ9jr�|*O�|&�������O�(#��BP�����vp&"W
�6Z�#R�#��,v�-�'9K�q+3�C�wz��!�'�������o.���s��c~�:R�:-�3����Gz����4M��'53�m�&gJ��Cc?P !s�LL��M�4�Jsy�">����^��:�=��pѵl�)�:7?��,3�����b O��d�:��*�A	(�6�?xB"񤦟��=)^+��U��,�O��L�]<���D,����l�R�]�.7�����e��*Rp�<I�d`�s�d�I�8���|	s�xTz�Z~ .���I �:�e��C��%���	���N@�&��S� 边��N�r�@��n̡���*�F~�1X�9~X�� ��]�W���L���9��?nw:�����$m�q,��݋�r������,<��8�`���ш�z-���oy?Hm�\�<8�G�����ځ����3�+�{=�� N����n�N�� ��^5W#���5,�N4��| '�f� 
����3J�N�����E��.��%�⧰�q�E�߫��-���S�$bo�����G)�١),���Ӂ�M�bz�fe��?_+C�~ѐG^1FR��Y>w;rv1(�B`ڢ��j�ߙ݊6�e�g�{��~{�zTWQ�����*�G������kn�vLicU�?��	���r�zq�~a��4�8��CsX�w:��hR�z�8��u��*%����cg�a�Ȼˈ�D���b:`E�ϓ���*���<k):�g�cA�8I��n<\w��֤V<��Z?r��v�oy2�~wo2�W*�<�ꛩߘ>+��{z|�R �[��;��m��,�c�x��A�7�g�|�)�a�5b��6�p_��;������kPlOT��ln�I�nU<n����������`��ڊ>�ەG�i/�x뤒�/{��b�	�
4�q����
wE
��I�tȦw懟��Г[[0�nk�+^� �=bc��jP�g��wѬ�	���]�H����*6�C�>|;�����������c,��l��f�Оj�)���B5|>�����V������X	�)Po��5�Tb:؋G4~;A�������dc���0r�?��*t�"�ZÛ��c@�Br�vߛJ��{
 K�O��u.2����#ι�7tΘ5�A���$�?�������)�Iy�P#EAv�	����u�;"� ��}'��,*���z��<7�����T�Y��K6K��e�PE�� @��WbZ����� ����
ģv��پfXϰ�v�������ez�j`�B�~Em��{@4�Gc���)�I�u��ZP݇T۬2;vPOy���n�@pUzw@	��̼&��h����Dރ�wv��^�=)�*�w���� W{���h^-���Z'-E�|>�.CZ���瞧�/��她3�<�ł7Jk���5g ��,o�za������`��ʛ:�4������ b�q��/,���@��یi�@�k�$�: ��l��R��~P@�x�Ik�/{�ˡWd=��P�s�5����оy�߾�Kʱ*���}D�e�x�"���e�nO\�{<}m�zOm53q�MQ�i��.~��݄
�-�~�=����1:(���U1-��7J��8� �C�qO�� �0��oJk1(�g�(*߹��˾W��N����!.��a$�c��I�*�n5�BV��3#p���4���"&DT�@�c����q��66Z��>����P4�=��p���@�SF+ƨ��M�L�1��_�ts0�7ԐSEn�B8��?�A@"�wLm�V�ؔ.!��#`��:̝��������}���_��ڃ����.̑ˋ���ĤO�O�r��S��i{��x$Y������>o��ҽ��l���m��uL2�z8.Uc�D�<.L�9�caVg�( OA+�/~���F>�^{c1���3>���Ը��P`��ǫ	]�j6�Ԝ�w��5���ݫss��z0��8M��LT�K�ۿi�߱�r��# :���Ƅ�v���>5�J�R_!��6h�0���h���X��|$��b*	�M��f�/3���6���U<n�F��R���u,I4$t��n�
7Lyԙ�3�"m󤷮H���,��R��@m1�o/U^�,|j>��"8*�
M��hsaǤ�d���pۂ#��/��X�v�9/	v�V�kߣ۽8�h&YC������=��w�M�X������O)�[W�k�����,��s�N�Zw��!B��
/���v�J�e��ƈ�!��%�b�fmJ�j��xE
����7�M�J#�
y�8�c�\:��(�����T8��lM�8
 ���qv���@<�S���8 ��7��7�[�f(d5p������ϧ��o���a>��OAPcZ���`+�P�f/����? .w�ߘu��}�佖�祡h/��g�?}~���q���!�X\���iv�����M{���� �d���k{�����
���
��kl�Р�x ^�WK�#��0�`Q�RM[�@00��0+�$����<:D�d��vlˑ��� �T��@^y��@����i����@^�����Pn�3�.[pS� � س���W�hۏ4T�n�������gp�A:3���(�������d�{����S���ỹ� F�%;��-7w8y^(�yV�����h	� �ΑK����a<��Ǹ� i��&Ĩ�����kl��d��8���_.8P�jY�9�Ϳ���?	hh�����-pa^$@��x PD�aU�]��;�N[��]%���
�tpF̽�y=Bv��A�Ї��w�����v�;��B��u������V<�GZ^='�Y�B���D���6� ��fS��d�1��4���M4��]���g.��9������HE!(b�L ���ߴ#3R$Q��;[���_݋�E ���ƤV%y�k?0�� I[��l����3*b�pkҞ��h2p]N<��ɿ��Y�ҽ��r��j�p/�k�"��"ܲApĀ/ۨ�kSJ9���o�����)[:Y|7�P��B�6   ����?߶�򛰵���E�J%��qb��~B�/Q� #p�4qo��jİ�8�F�1XwOe���z8��w�̳��h^�^�S6y��C�2�
���&+P�Ȟ��K]�.�U�fT��"����0MlCޫS9aX%0df����`���6%�:X�B�lO]�ƅ9uo�">%��T�ȼK������Fm&���S��7��E5�/3��[��:��c�/�`���/��w��L)r.:%�V|�n�����z���������mt�^���L`�	*il�
q�n��Y��nĐ��xc3��J���n��b5
H��'ɛ �Oype���%�,Q�J�X��R������5��6�TÃX2��?�����R	�d3H/�^�S6*1�K|�}h�vԭ�R��c�7~�9���Ak\�n���>{���m�Y¾u��.mB����]LyL˨w\��?�[w��/����v/���`��"�d�ҥ�P�����e����q�?��0̠?�[��E�1�p��@��]��K�w���.t�f�&IoK����g"�+[V��5�����<t�y4�d�3�b�����uK[7~���k��g�2�����:������w�5� ��G����������������_c^3� ��J�y������_��E�ڛ���6��C��%�O|<�oז��r���,�?�aO���6֤�˒]�s�C���4�(�ZG/&���X�:�f���-
3-�R�I�W71���v5j7��਑Þ���C'.�B^m7yl��{�˵?�n���,�����9�ܽ[�s(�ȏ�<�Kcm�I���xfs�~����~Y��;���c����.�E[���(��6���y�3Pcs�#rq���d�0u^�B�����}�����7�T��p���W9��>�P�W#�R��af�o�,� vDxs�waQwi��o�ǎ�m^Ӿ4<�D�{�9�U�N�ouj�sɲ�VR9���ț�6����(K+�e8e��k�7��n�3��BԯJ�����87�x��D@�޳=AAqHG="��ȏ����uQ����D��d"}�^�cs��n��)�:� �%ϴ�:�T�4=�4t5�ƶ��|���|�g��w�nZ4H�s�^�2!��O�<ʑ0�ԭ8��-��iz���mw����^#�;�x��,/}��qm3�����j�!�_jD�߅Eg�SS��jc���jsH�ѹ�Q�X4��b[0��#�?D�&�of��KM]��G1;~���s�~Y�a���
�^>q��;��84v���z6��3��=���59=M�72���h=��j�9B��&~wM��U�K	���ٵ*�g�W��v����V����̬Y|��7�.�vQ�'˄���G֙EJ���?�L͐]��^@�+���;<7��a���E�2��w~"�c%����ˌV׺\P�((��'�r�Z��b�l�߇q���qo�oq%�#��=S��2��v3�J�A�!��*��"��q�k�ʬ��~#���<q6�@ڙ� w�ԁۖ�{h0{Ű���(Y���oRE���;[zyG�z�7�v�d������p�-�:m�҉иk�?U}׌�D@n4!���Tz]+
��H���M�d��u��J�E���p��i�_Z7�9(�9�S���l@���Y�ny&3,�-aZ9����[��p?�y�,v���g��(E�%�?��k�+������|W+!�|x �5�N��'����ŕb��Q��B�.U�]�2�������7�!6D���9W����lH��j��Z9�F*z�85#ńH�(��4��?��ѽV�zJ�k�
۷��*|KU:-�D��B��|��u�m�󙀳 u�,9�9Z0��U��M���R��%�&4� �	ŝ�|�<��*���:�ۼܑIs��p
r(�ĸ�몜�mb�W~f��>�/e���A55�$��¥v�x?Af^�j�Q:lKD�XR���V<ݿ��BP��tQf��a�J�����m���
5�ʖ6��I��BJ�Ⱦ���R�P	�P)ʞ}�[��k�dwqm�~���]���<O��<�{��|���y����o�6�6ba�.9���&����e���0�Z$��3��je;k6�Kl��X�?����55�ܥ�«'��Kf�r,W��N�i���ͷ&��k���L\�����7���ǲP��?y���4�0�D;���y�+�#�����ƫD�:�X����������Y4F�Q�J(��;�j�����M��-��:y��qb�a�H{߿�o$�+�KzM�-QtM��w��n�Ƥ�5��UD}ll�b.�Ո����kRZ��P,�2��L�sơM��U,��D{�� s-�h�;��Y�c�H�"���bQ��;�,��j7�5ʻ�]�w;�/k��wTM�L�s��zl
��t������] �K�S}��_T|��ܓؗ�1�dd���?�=��Mm��ء�T��5�(	�Y�@�i �;S�_ؚ�!CT���Ua��&���°��:���S�h�Yev��J�Vx_Ul��S�!�Ff�vOms���4�ԧ�Ш�9�a��xZ�X�H�s���f����1S�cv��&ʁ���	Ղ�>�Eɬ$b��U1��&w�R|���n�$ߪ����`߄�C�� l��&��V0p��2-f�|A�W3������+Y���J���Ҋ�.5��=<aLq:�v�Z�&u�~`n>�i���Ǆ�NF���XV@}�����j��)R��U�ַ�Z(�r�}�@Ǽ(_�x����)�\�}�6
K�/�:M��p���L[�H�C ��oQ�`N�V��\�᳀/AL���wiX�\��V�W����"L�S@KF[�\ �%"����/xQ�^�$ `~�����L��<M-�HqMUZa�������V��\�k����u}=DQ����~
B���i�A�9�����b��c^�	C��l�VӍ�t��rW�8�~�2���]��d�>k8���]�6#��YHu��t����^���:9c�F�^ڤ _�����hN�Q�uu�h�����¡�R;\�2mc3�F߆���4�yg��H������s��<�,P�����W��*G8�Ԅo�ų���"O*��e����eq��KDԈb~8w�kF1{��;/�X|q�әj
?�����`m�@@0���3�7��3�	�b�����_��������?3x�1����ѻQ@Z�(H&�Kз��M�n��1�����|�L�˃E�8������!'z5ج#~H�w���M)�u7�7C����[�'o�����uFSs_�`jX�d"
��P)񒶷��///@d�Vb
��	ӌV��`�xn\�^�C�<n���t�8�4�N��Y�:�W�Au��ڝ�]�R��)�jX��sFU5ܔ�W��Z@�IĹ�Cq�\o�����qV\�܆z(�9ځZ9��*�c�.G[����`��'��F59�A�Bt�����k����fYi�޹��o ��U~4#-�N䣘�R�͊Z�,�8�HG�P���B�,~�V�*A-�S��و�4Gr��o+�~��v>���%p:���[����~I�VB��y���Ft�F��A�L����#���l������zR&i��+�O�����@\6Х�xO�ʠ�"����pK�6/�0S�r�罺§w2Z��k�n��!N�u�x�W��(�W&�������6��P�t��f��<�����L�����z�<�8�JX�\�[��;���쮓t�s�U�4}L���o�pܿ1��Y���[�FF~�x��4�6.�l�������x����Jt�v�T�p'R�@\��g�@�x��f���z�F��y��A�1���;�j�%c���v~�����{�~�M�YOR��S��Z�	#\�"����rfh�}�hj�i`��oR��6�Eʸ�"1�ҹ[s96���$��OZ~Xx���I+�p��;��V��g �`WT+E�b����^���Fr&VH�*���|$��b�I�~JPw�#e��Rh�\OT\܁��B�11�j|��1s�rWtտ����>@��Hpz9�i���U>��e��dĽ 	NT�fƛN0a�ʵ�j���c�fO_(з:�$F0n�*o!:5!�g�t�%_�[�ZLe�ۥ�c�rϟA}���-�5��/�)��1ȟ�rkc��V?v
��+%�G���H���&��(d� H�F-���[ǜZ+��YX"T ��₳ ���D����!4��K~�LA�3lf��$&n�gd��k��,V`B�������LOv�1�uL/1q~g�V��yP֣�������G�� N�X�Q�c��@K1��+�A�-O�U8Pر����y0`:)~��d��N�>��fe��k���FQ#VyȂ��T�VP��ll]�!���u���#��x�Z�fy�)D����eȮ�a?6Y�r�.4���C�iὂX�R���?���("?�~���S�.G$��o��y���f�5����:3SZ'ԩ��פ�b��6h[�ܶ��3�f��At6��(u�k�� rg�.i��E�t%�ƍ꜑�T.��>�H��s`�)�En��tN��Fu�=4'��8��*��4���\�>��'�y,����F�����Te�y$G$6�=��H!̈́� �˜�൘����e/4���jZ.��˅p�����+T��bўˡPM���N���yw�����
Uq�q�wW��C����ܿ����#�Ν��@���h�񕩪\�D��
��eo\ܙ��Ƣ��

�6�b[Or������I9�6�@�@�����@�"�7Q�y6AVAf�ys�㞹.i>�;`�(�q�ڍRMd\ʀܨ�2�VV�Ke�����SK��{�S�����d		�ƙsx�鴇��-�ɼw
�*z]�}����Ź�a
��kp[��?�Pe2r���Y�
��f/�!�z1��S��PX�Aisb7����?j�z�Ĺ�@�,cCn��׹�������`���Mqǟ|"����f�����2�g��^�s�������b��/��M���8C�- �̯���Seݮ�?���?B�}�_��{��8���  �����6Y��ŭ�Q�5����\� lg��t^��L��$�)�|��:�fj@wVBWd`�g��U�hn��(�R���� .gR%��Q�O��d�~�����`?�ȥ��b��%�tDN�\�dOߞ����ƙ��ȓ�����������:����"%�ڢn��I�'�F�.w䴆_������\�����7�G�#C~��fr�J�:��u�m��{?<e��jG���~�vm[�zltA�X:��j�s�nW�Fr���mɴ#}�ewI�k>�a�ϻ�ϿGn������Ѓ�;��K�^c�I1�G��h
,%�k��\������( �le��\S��ڭ�'X�����&�2��%�FY�br7�|�;���L��v�p�&��#�'��Lk�O�Py����;z4bXd[��̞�����+9w���TJ��'�1���Rp9�:�6��[rw�?��G~�W�W��?Ż!FԀ��R�L�\��Izy*�ea`�)�t�kBN�^69�a��Q�n5m��skc�45�R�n8�ޣ�?�B�3�G	���$:Ɲ��e�Vm��'g�<'�^�>���ѷ���9E]ޢ"�[��ߠ|]	�-sɥ9��$�ǫ��4��3m�R�'F�'�:կ�4dw�|���[���P�)�T�CJ�]���#��[�k�C���9�����	Gth���:�s�Ĳ�����XWԃ<V{����ϣeiN�af�w�\D��������yH�� V钰>�C\��� �Y(�Ny�@�9�XE��3�x m@z���&�"��]�Y0�p�c89�\���Ε�O|�*^�Oy��x�a�l�	���i�S�{A� ��������3o�)#d}�\�r��#�Ȭm�W�vPf3�A�	��0\�G�������Ƈˡ����Y��S��n�_��[�d�jy`u�s��3SN4�y�Z`��R]a����|���xJD�{R�/���1/�*`�1�����lk���5�yxo%�tU�� �S������3��FHص���h� c'y��������ӌ=MPl�;i�5V8)�#|�"�떳���{h��;�v��bg���� t��,�K�B���ˌK�Z�R���܇%��Ʌ�:��M�U��&�!�"���ܐ���U���_.�--T���ڙ��,�������/|A�kתr���l���>�����̛�S|���©"&�(�:�xK��D��iHH���R��n��a�=]�����_>��j�����>,����U��|�{���x���O����t�:ک�\����	{���� ��>c-E�qc��}�������KߊƇ������IqI��V��V�s�2���߸�s��Fw���jIMߏ�s�Cj��������*�[K�[Ϗ\��+We����~�ii?�,^�s�БQ*����`y��i��|���k�v�C�iw��3�o����:7�Td��q���5��}L�.A%���<��\��������:�˻17�=��A�(���"APuߠ�����4@N��UQذf��f��S]6�y_S�a���"9J]��Sk��*\�Ȧ�WO3�awid�hR)���L����t���Ɖљ��<���������B�!19�L���ʬA'/�cx�{���j^{{�!a����
볖�)#����W�Nc_�R�W���a�A:b�̐oκ�k���A���[ŘR�`��s��l�֢��"�q��Xg,� "�-�,�&�e�2P̡�o���8�9K�e-������ľ>� dЌ��]z�5��ؐ��!�7��\ʫ
�0q�[^|ѻ@$��}+�ڧI�;'�A'�O)F<����_�~�T4_)E��M��>~���0l�L_��pu��9C~�����Gy���\����ƭ{X+ٔX�@���K��,��Wb;a9W�NhK����*���'�;b�2&��_R�.'ks2r�56�˫�;�5#��G~w�֡6�B2������x�
�ƒW�=�b7�ڽ�J[�5H���&���(5����>?�4Vh����{rO��d5I-K[��ܟֲM�7������YS�A�Aw�+
o�֚j�na���{|��}�6�0���&��d�d��q���CaQ�~��Q	Uf��4D���{vŠ o�1�'
i&�.cQ��n��t�o�ʉ�O���(���ɫ�63�4*/����~�f��%bS�J�Hj��{4��v�Q������T��C�Z����Vz��0��-��P{�֥�%����y�*���j����ZOk��~����jk�А�ֈj�(@���xv���H�"�ܙ �=��)"_1�,���q�ڼ[�|kA�\c��]�˃��_����;*�z06zȓ��<����WŶ� �Q��3q��$�r�M'Yo�VQk7�zSsF������\�'̗`����_M:RY������n|s��W1Nt]��4�K �)�i�*������'V�#x�b:P��������	M���P-;|�|�j���lF#�>��}�N��iY��%+�/bpsG���w��i���d^�v���Y��	Z*Nr��~<��D�^5|�e���P��'XN�[w�{�>g���jp�*�DG&*�N��!�����z��	T\vm����c׭ڼ��|�� �zR��0��I�`6�y·1�����3���Ip��7��`
���q����~���r�����X5�g��9k�ņ���o>]�Ҫ1�3��gY�n�"�19��6��F��*'�_�>oR��%�K?�yY\Ԭ̝i8Ծ�OcP���}�W��m#������|����T�����Y�R����wc|j���zF%�J��;NNUe	<��L_�$l-�a�iy.T�H��Խ�N��]z(!y,]�1�WeP��pV��>ڕT�١�HG�hܦ]
�nƒ`�	t�\/�,�)��l��W����%E�c)�E��h\S�k�a���̛��Z��Z�xd3�P�mq���Nr��Nc�A�c˱�,�VJW���9w��@ޤJ+�]j�Y~�R�㢟��C��9(�!I�_<å��p��3+ߣ�!���q�H*Z��jM	�h0g�%"*�(͉�$R�s�V��{#^��^N��G�r��~�\��3b?ΨKw���HmH~u��U���5�5�O.r�]������,E⨜��g�,�%�!�ʺ'�+�pn�×h�D�w,PںI��<���H|c�%[3J�|;�����\gnR	vJ����V�H
�6#þ��GoU����"\'���S��z"���q�<܋��T8���`�EzHQn6�:&��C�͖lǆ��O��ݪ�����y�l���W�-�޲�دrq����?Bf�0���S?��P��9�tD�8�}��%���q�s9j�dɃ�[�X�������P݄��.�D��EYM;��3��ѽ8���#�����Y�PJT{�x3�+v7JJ�����;��5���g�4����a~���%=@朗,u�w����1�MWŮ���ѕj	��
ot�>
eDޠ��>���-�����\i�}X�hWoIR����4�H��L㋏�Pa��3�r���7y�0�G������2���#%�����*�3��ɪ,�n�H>��[���1���El���������R��Xy��":n���oo�wN�\����[�?E�xO�ڛ�-�פ�W�D�MԟmQy�3pf�>/�l�A�x�g(�cz6}�2��t�CQ�� ��VE/��D$��dGN.��z3b��Y֒V�Y/�?�����Q�t'���Q2�\�
戤/�x�'�E����;��q��G���1.���9C�Zu܃,�W#��䯏wU�w�����mZ�
�be���O�i��{�&k�\�9hK��y�S�X�&����8)�<!�/h��x:���#V���nbuZd��|
N�E�8�u�N��ب@�xs��G5�Q��{/�b���r+"��;����8`�\�M���'����4E��hSo��o��{9>�-@�x�P̳��1�S�^2i��,'�[0e9O��cյ��ɾ�T�݁��(�-�����4p����5¬�nH�䙗F�e\�Ëw��Ji��������3�u�&[z.�VX|�m�;2�pN��&bH=�)�}�^������5Jj��2S�ac^��Ɩ>���?	g��C3�A{�5�)=�F�5Cب&��V������D�L9��k��4��=<Y��Ҵ�)G��)u x��ވ��>��.C�L��!�4b��7�Du+-� �������(�<^�h���wu��?e�v:��|����v��>S܅~�O�7����/ѕ|ƺ�;���L,w�z�M���D{��]Z�i.�J͡�������x�}E�Bk4;G��ڏ�ʁ_@��'�4sRyNM�u/�2hAـ�[���e�Zλ���}l�e0W�nc�WY�@ [�9)7\ɜ���ʊ��K�ca0C�E3$8)g�Kb�K�$�h=]n�=(�<�1~$�u���}5����u�ʽ�BAW�t�8[*�k��I�ً�Y�����R��rƸqo�s��ƌ�.l��KP��KާB�����^UCN�E�)�rhE�u~������TM;�`Ne$��>*2 ��k.E�E�8Xd>�7��ZaS_�M�ٿw"�B)M���k?HL�yW ��*�5��D�L�|l&���N"Pj.M5���2�X;���y��M��Y���Hޑ���c���j!�Ŋ6	�2;Fms����RA���<$�/>���r��ċ��H�r��dXT#���+2�9&�+~�c�0RJu+(sX������a���J������O^��n�W9�l���ف��w�_�tA��Tn��_�m�x������#���>��[���y�i�v�Gh�+u[�>V"r���4(���q5IMVYs�%b��`Y��r�;vX>���V��dx��`K<��k쟟S�s�Wþ�3� �Hf@O��Vw��U�-:����)�=���c@?��Ar����n���f�pN���]	��M�cfr'ܮ_3�5-�U;�;��G�2n�Ug^��䶴�/	KX6D4��_p2�s�C���H�J1�����y+��I��~�H�ے_Uu��*D }柿	�C�w�� c�̜A϶b:4("a�{haU��B�C��ϵە�h��:+���;��@FB�����G���]�a�(�����vҼ׊F������?�Y����ӥ;��ɍtNZIN	���#S�C�V)�B�O|6֏���E��U}�'�rx��ǞO�Q�;��u`]�zvu�E�p-��������;V�׊nbM}@S9j�,#��V��Y��:vGMџK#}3��b쐨D��b�u� �ʣ�!�l��w(v
^��QH�����=yKV�� \�I���Q�� 	,��I�7SX�Kg��n��Qуd�����R.=�V&�u�:	9}+����!_6\Q�cݘ�O�Z�����b#��b}�\n��t��L�帋>5�ƴ��p!�5��*��䰺#�T��`�2�<�b����1�s�-|v2�6ND?g
/6��"�h+O���e��˒��ZQ���-3?�9j�ʑa����1���G[�`�m%M����X��=�s�nNy�����v[��z[��*��T�����lE�T~��;�KP��%r~}��%t
 䃆��!n`���Vڤ��r�י���; ����ٲ����-N�F�\s�I� !D���;�'�0���W��$�6�vG���
��I��P������+�o&����N~؉Uў�?
'�,&��V
!xՔ�'\�dU���X���XƱ��� d�6֠�X*�E;1�R�[R��ȹ�g��f�![���]�D�����εl¿�1�x�X|NQ���꟧��-M�!>L�?�|?2\��G���L��k�f����;~ћ�K�I������^e-$nWv��m�鶵q_�P�����'e�<�I�.;eǎ�-{C�܋H-����e[�-�Y?�	��v��su�����ׯ����Mc//�䱗32�D�>]��á1�h����H����G�b��5X�3,Y�=X�/����Q�Kf�0ӭ��e����W"��z�ܟ���Ũ�I��p�����1�t&j)��^��E�(^����ެ=w�G�=�i*��R��-��E��}���G)-G��l�B���<6�x�����~U8��C�pv����S�K����`������--1�.�K��1�gPfa�V�����53= 7H����)vO�sd��I]l�k���k5�s�%�w�t9�B���Y�[��l1����ɞk��ac��^n�A����7h�blV�/���b�V�?��>2\8�]��Q	Z�s�Myj�ި���b�D�5�Ǘ�����n1����$9/�q-��w^z���Arx�����ݳ��Z��	Q���R�q�z�"Ӹ���h�HwU�E�?=Ό�;{����K��:Wáq��F�L~ɒڥJm#�����s��|����࿨r�ԝ�e���
1��z�uQ��{n
m��,{�fyF�d�r���1�0?�����]��EX0O]��{K�x�ci_)�⺱���k�,f7d$Jԭ�����g�J�D��&K��nرn��8G�Q�M�u�>�2� ��S�e��ײ��X��]�:�?,F���N�/H�xL,i�١��i��ҽ��L�53��]�бīt��T֐�����̏~U�Ut�������=��}�{g�p"M�t1�D1��W]_�?Q��O�/�R���L�nmٕt�p�*�Rf�JT,���� !��e�0����e����cӺ^m�3+���?me�*��+N���? �e�1S]#c���ެ]���d�K���Xb�Y�^�oWr�x��쾞zeކ�����`��R�j�����e��J��i"�T�v+���%�-K��OmȬ���q��䑒�-J�����ǘ#y��ړ�9(���a�Up��.G�L�.��h7X<C&���11z�މ�߇e��?\�^|�l�Ē�,�%.���G�\�X>�l���1�ǃ�ڄ�>C�G�6�z|��hG��<���_��U���e���B��dk�B)���YY;����VpEO�:ñk+�[����FO��'D�<�wk�"��]�ٟ�1@L߇n�̜��qv�p�55�@�Gߓ�	aPKC]̊�3l�Y~�o�3^o��T�ڔ~I�T~lm��T����xM]Y�d3��w���n��.l���/���8vo�o��)�~q���"
O�6�=�h��|������Q��ީ-�i��p���zv������F���npa�Д��%����w�����-G8��BT�1rz)�@6^����՜T, h�u�*R.��ͯ����A�i�n� ���.}���6��;�dY��4d%Ir��7����t�/�]f�����z���-��?�|��z�2y.��wh�]ea�"]䬭�����$�I���c��ĳ��ʭ���u�7U����1f��W�V�x�DA�Vo�,ߝf����O��7c�뼄��o<�=O�;�\��K�>I���A#!a9��SC֮��ȇ�����tؼ��EP��
��nj�+;R����H^ogo|�4�A��x�ɬ��R�&_Z�쫳��������H�}a�ʚR��"�t�ȇ~ZG]E�ԟ	K�����s�ȑ��"�Y*�[\�UHF�"X���j���A�R�,X��3�q���*ƒ�p���U*E�y^�$੩�A;�s�;Ѯ~h�y7j��� S3!6s�
��M}�c��Qʺ/݌|p"���fT+����9<&@��*�Ƣi�l��`�w7Z�(�C�{Gl^����H�%��c�>{�׎)'��!Ə��N:%�s�;W��63}|f 8y$�F��X�%i��m�j�xo��+MG]N;N�eo���Q�����!x������ʦoK��ܡ =%��a���;:��ۿut�������'��q{��;����*(�:t�W俘��q>�??g��h�=?�&c�P�$�w�,�Y�S�Te�zr�*ƥEa�8��}*���u`�m�I=�g�n=�1��p�OW������k3���O�#f`.R��h���n��紼�L��>M��|Zs�nތ�%�����57��c4�R^ 3��9
���37��oEmL�!�^�(�tQ���!�E�#
$���]w���N��V/z���,~-��j�� ���ͣ� g�͔̈qD�nQ����á�Mj���j@�.{�EL@mм!�1EY�MS&"G5�����85���tՋ�¨I�	
�پ/�o����9YǴ�r��5�{U��>�H����1v�-('���o�aKs�`��`�E��r���m���t���[��ln��)��nW�#c�Ò�Egѵp{�ô��ؒ�-��zܢ��'@O+�Ǐ�����TmEAe���n�L����w�>��s�����G�\!t������>�!��ѓAU"���[f�*�Kq4���1M���,J(o#���E���eǦ�)�8O+g�G�OSs��Oj�,iG��x��ސ���૟֓de�OY��>dc�2�bÕn�U�tȊ�Y?����8!��>M2�_����K^�{����I����Ȥ�FW9Էױ!C4ҷ�,u84��u)���}�[
6a���{��vq�����)əmb��}��r�ec�HQÖ����&�ǅ�|�4X�:]�"��p����i�<��U���lA4��p�Jb���2IE�
wT}�N�(NcmgP�Y���o�(0��0�Ø�|岥�=�=�|��=2�xf���{:�����C݉�g��RM����yG㝨ޅ��ɼ,�~8��	����9A���"��ݼ�@L�!���˝�}�}̑���hɼ�	�`g/Q�+�0�N�<��Q��m���{�|4j�
���l<ґ�!�yd�>�_xR�۞����,�,Ag������&HB6��V����IGbo��gz�l��� UXp�V 丹��cp`4�E�͋�
>����`��5���6���<��>@�@�L��
��[/$�l�Ó$�5l����䵠�[�,�3� 뙷n񖎋����C^�4u5ZR6*�����?�B�@ �.���_����H����N��w羨�bb����K���O.^8�����p#F�]�J���""�P��꬗�Q��Bv|��1(j�R�dM����!�\����&��|�H1I��X�ՆЙQ���K�
m�L��`��Q��V*��0���K0��Dex�XCM4E��r���J2��n�{��K����1[Ϳ��哆��M���b،f#�6"9��.�Ab3�K[b�d>�?uG�=6��:����Э��v�U����NI˶� O�ݱr>�O�f8y[�ЀL���c��T5�g�W�Xo���[p'� ���&��r|8e��,�߱�� J���Z�j\Q<@d�8����ӷ��"�߰����h��j���Jl��˘��}V��S��8�`vRu�L"f��_� %d�%Ǘ�+�[��r�����?;:��4GE�:'��_����O3��ġ�	�\`��[a�ۖ�R��� ����u���&�0ҁadpI�WZ��VڣfM��d �䥰����I	��mx�1/�����G=�"jp��`� ���Qu��U�W��)f�����а��ݻ��5W�A����ڪ(��C��+���4|b���TϞ@'��$�`X]
��--ݝhg�v�����VS�IW�Z�w���V�:�ڋ��}
b��	a�Ӿ��.\�I�q�t�`?l 7|�&n{��U~QF��*���&[�,r������=��]Wj ksw��`�y�a��3�9�b;Yf;� ���O�	���1��W{F) �g2m�� Lm`m(�ci�=z����Uzz��<��?��䄚�Q�s�B��,���n馘�{./��[l���u�є���d/�KN+�46��jW�*6�rM�^���x�5z�bG|{�����`ׇ9aǜ�G]��Ū�Y}�.��6#�VSo�� �#��M��r�I;}A=�Q��0v����I([�����A�k�hVD���]��1{k���M�:}����lR�y���AA�u��=�H�����,(b�̺ӊ�r͞6G�(����A]�o7�n�b̺�e_�5�7�I���;��#��!�-Q�ަ������(�{�6C~��m���XdS�\*�	ˏ�(L���_Rs�\@}��`X7e�/��Z�p�yшF	T�HП�d0!Wk��q��P���! ��M�����	Eb�57E�����f�[X1j������&�PY�{ڰT��Su�䞇N�c0��6��>��l�f���L��a��@����N�#{�v��[!8���*�;�DΕ4�hU�E|�C�T2ѻ4V7�=��°�Ǝ�)S�d��G�GЄ�Xs
\mƭz�%I���g7�~9�܉O���-	`>����h�	��:+1Ú�@R��I Q~��?�~Is��e���;�ݥU\��9��F�A���E^�.�W�$�[�¿��2r~�J�;�?�:!��	A������&G�Qx�EIZ.)���`/&خa��YE�r���&���eW�7 .�� p�� �@�t2�n�fy��+e�«;
u7��$aW��p���BMzo�K]����g��T"�P(v~�z0Mw'��l��o�!�X�;~"\;�N=)�+)�#�s���2��<�*!����Y��f����T�!04�{J�`,i�����B'��uL�@���~f�L!��&Ͷ{x]����-Zs`���l+�
9X^��5�\��$���?�Qo/
�] �q%WuM����~eG�^�f��U�T��qƑ2%w�ى�J��tw.�ůK�]�#E�-�c3/�E���9U��̫�L������|��"P���B����ECڜ�#�N**�l�T{M�D �"�U��j��m�$::���~�NA��ċƨ��g_^�|�\��Rۿ��9��#�2Z	!��^M/Q�Q#��dz��n��f��� �%�)Pv�F�Xj��d�O�b;c+��0�ՠ��ler�ho��*����#S/`����C<KG��Xg�`�#��ЮW^Z~��=��6Z��{���Ŷ��2W`ji�ԵLWյ���(.��ۘ���h�`^�׎�~��7߉��\�"&Ѕ��׀���x5���WM�ךLAޡO�[�[E�/[�cjV�.Bf�6Zp5-T�̔�""���w��8�Z�E��a|�*t���v%�|�v��I��z�
�،�'�*�EO#�<��78���{�Vr��7t@�F�\`�Z�_TE0@�i��w��/�
��B���2&|a��ŧ����W(�NY6;µ�R�a�8��('�#a��ՂH���� rd�$�2�m`�E!��r�%�6�})�|_��;�
��'�[�#�!d�~��R��\C8ƺ*�~��`߹~��6��W�
r��&�;�Ծ�\w����/�g|����K�ĳ���~��t�ɉV���/��=����@q����v�������i3�w[�o��-M����5-h_����3:���p̴����i��ϥv�XT'� �h?��x���W���p�k7Z�I��4lc!�X��x3%�-��Q�Հ`�F���������@��_����l��By�]i�a�=iF���,�h[�*�D|#,��y����̍?���dV�ykߍ�	6��b8���A�?7Zl��$C�������>8]�g`��}4~�}V�R�K@{�k�TT�?77Є �6�fʲl�.�@mxSr�Q�xIL�Ƅ��M'�/}�r����X��r��iR'C�6R�sP;�aÇ�>� �0�{��P;� X���&8�E �F�n2�蒱��:L��@��u��Ƭ�:��������v�?������F�`�N��)�f�<N�)[5(��ϟQ�~	�"�f�(�V�-�!�۲�c�+Ńl�M
n��➻�taq�P	Ƿ�@C%�moڠ�t��U
R޵�.��{�t��&V��;�G=���n��Kͣ,i�k�YIM�'s���R�{A�V�k�H�T��~r���&T��"���%0̴ ϥ�zݫ���x&b�碦v��~�Y$Q}4�v@�q��ǃ�-o�����<�P]��ź�`'k]���A�!��D+�]x[������;<����OM�'�3c��ı����Cs��h����ǟܹ7XȓrX2	��,���%� .*�q8����� :uO����0R,�;�����LN�6�OpĶ����>��2��˝�tKf�:Bg��{��J�T?͉�Q������S������0���C4�
�Cc�7�y	��#�{Ba����/��x��+���k�Fy/i�`����y�DE�A�1+�mBG�������+�|��H�R��-w��.�u��?���B�YD�/�S��ʜ��L�{^����3T�?�/�.GI4wd���ೲ2HB���4�/�ލ�����%Y��Gɀ��2x��7T�Zi�s�p(�A*M��0
�n1<5"�㴥q�� ��)1��]>{��$ġ��5���o ��<d�?ZD�z�aDz�i=�6���?R���4�Z7�`R�z�z��:-"����}p�3
�������i%xe�E8�A��/6Σ�-�_�������ǟ!˟ݩ:�l��Ʒ�]�N�ѭ��\[UN-���
H�W���_��֟Ӱ��K�`��0n;��k	��oCT���X&��[=.�<��������$�zal둂-�^�
3�2�mē����O��a�v�T�ኘ���v�?^���o%`j{��Q;�r~!X����MҚ�!^��x_��A��m�?��~���-�p�3����N��)���C5�I����-����a2m���_J_�v�m��p_����K^����͟;���Rλ��T��ol�uc���S�ߔl/��V���'%�cMsCu5�.Q�3�W��$Q�8S������մ}��T����߆Ҍ����y9������=�7=�n�*>�lC��6�۸�6;��;���-��޷�bY6���Uߖ���H����0�'4��#�W4�R��r�f'�_6x�����t͍4���E�zd&�zتɼ�WB�G��}C���Ux{��K���9��V�#i	�3�
�=�YV����َ�$�{�3�-���
g�kG�o���Ic���	��&�8�g�����xF��R�2d�˦���XW>v�?S����TZb ʟ5��q?��m&x)Ӎ��9�Yκ�E��Mv��7�+�� GP�܎x����ʫ�cw�.�2��&�7��+�g�<�h'm�w�8Qb�S�ė�g��(��p4���zd�a����=O�f�C��L̙f:/$U6���������D��_��O�zw���
��H�9�>�'.��Ĩ�A]�y؍ʕ�|��ɒ�Z[��(|{������ξ�����#�ʡ~��[�g��K�ۚT�t;�eKY)f��yN�}�c�B�?��2��K0o~D�y���Ҏ��-�z&kx�"�2�o(�n�$��ܻy��=Lz��w�??Q�U�~�j��[�E������-���f]x)�}Ӗ����@������'"2�û�4�3�����XbO���[ҭ�\HԽ.Xm�}��07���T�~��k>\0�����?[ұ��<���*9f��L�ts6O��<W���~~�e5�M�L�0'�'��ue_�m±'���{�+�FZm��\]i $�6e��x��sgG��58���g>�� �^��w��>�
F�����b�0]��:�:�:�O��ι���Bp��֙���@e��f��Χj+ l��g��,�	�q��)<Q�#}Z4 b�K�2���nb�r�gs<[���������3Y'�-�*�pG3W���=�7���`C7wu���\X�YR��e��$��p器ù�&):�8�iQ�&������z1���k�	�ҕO��t?��� �[Q���m��������=���E���:z;jEe8����[/�G2��,D���7=��q�rp����l k���U��d(p<V�������ժb��X�C�\�i��B�KiGfs�C��@<^��bϒ��7|(bS�zq��UE��k��@�8�Ù1g��<� �ZyU_�V�V����P��b�zp�����h·���n[�M���)����$�qbh�r�y���DW�G�N��u��N:|����4TK3AP�dxV�GQ
v8C_9~���a�L+��N@%)�%<}��%�ֆ�5�yBz�wo�[y�IEa��4c0]����v{!��ldĸG�7"�lL��i�Е�����8�ȉ��6�m�� ��J8�>��')n�%�����r�c�:b��<�^�}�R�#]�ie�I��HGIԽ�� ��+��	w<�,|L#�[=��������K�S�L�S��qEd��7��ᛧ	���gx����1�Q`�u&�Vփ�I?GͿ�2�}��7:	�"A����h��BH���A_�<g�ee���>������;�(К	b���1�p���XKn[�F�S�{���_�?z���8V���H�zQB�;�� }hf��{x�t�鵛C�{:[;��@��Ղ�)=�G�#
e�'�{ծn�=�;�d����pt�'��>���l�8�4�p0Eܜ�b�c�����g�/����eY�g�����wW}�Y��]��;A���C� ��˧.�.wJt銔u�T��2��B`�����؟���k{�ڢ�ޥَ������eVb�w�����)�/�O�5��?�z�"�W������{	��=���?�x�1��(��TZJ�V7�v���M�O������K�i�rs�9�m�>	�̟�����&���S:	)�e�I
��iяmeO�Μ�><�'u��ڊ�=�Y������r�F� ^�*������>P[b��2�
�<F�'R*��C��s~t؊Z�&'������Vҥb~� ����9s�#x'�_����\�-��@\�W�k��9�D��j@G��VkĐЋ��~�Y��v�����6-��8o�����Ȟ8��	m�Ԗ��_�0"-O7/�}��6�g�"�4b/]�0>q.�RT��D��ƿa/J<�vQm��%�<�g B���������GB��ľ�ס�]q��������g��eM]�v���~:r��{Yw��4/I6�^�z�g~!�W��[�w��`��>����r�Y�z������>��p��1�'M��eyʊƶ�A2���R_����_	��P|�S��љ�C"��R�B��$�3���\��ů3�.N�=|�T+FAd�B�6Xj<c�����5����{g��D���@�K�mpeM�g��W�< _�+�JT�u����/���lbn�m����}���n����g�m�����w����)���i���"��B'�Nԫ����WY|P�'�i��'t���w�sp�bh*�,�2h&��n�$4��=�ljm��( "es����^�]ׇx٨9� �/: �q�#�?I��f9]���ȎK�%��",�A�d�5qH���/�E"�E3`�]�)k:k
��l<q�ϫ����.�,,M�{��6B��#�yl���>�M�>�*�HG��ͷ�͑v�d
�/4���ׅ}C©O)��R���/h��/��^P�Y����f�W��F`�$�z1�:b�ˤ�s�ٿ���VÒ�9��b��k���_;���ہ*�
���*\*q��uRz$ބ��:�6_�}W�f���f�g��:�g��I7��{	E�Űj�ֹ��g"2����!ߜ�Q����k����S���	{�菸�����~�|�<�u���r1Č������Q|�7?������Ū]���m��3bg����-���9�lBBa�������=�ePq&A�߆1@�FPG�[�G��&|9�J?�&(2�h;�/�����޵�hO�f(���������G�&i����A�>�OD�+QVd\+�q�T�L�%{fo��yCƥ2B�#��<�9���_�y�����~���sι[{�i�7l�R���m6V���Ϝ������ąH=磨����T�c8G�A�X��LcsS��Sr��1��{���Dt�A,��u]k�ZW���;a�ᔃ߫��˘ā�T�?0K��$�������ˊWeL!�@b�u����T|���хI����1��ar탯{J�B��+����H����Y͙t���h�U	�oŨV�*�0��YM
����S˥Bw`��~�-4PUq]z�@)�7s�S`�p!�,c�Ѩ�c=�+�y��P��Wa���i�@lxj>��)ej�}x�7hQ�lNP��qQ��R��y�%�Tp��Nvs�m���bV@�i�<U�L�][O�'J�RM�����),��5ǅA9��*���ٚ�>U^5�����O�I,�5A�����1�#F�����n���:�@�t�tIfF����31;�9�0M�_�:,Z��v�n��_ �wHXn��	Y�%�0e4�-gݖ��4�A�ᾆ�ؤ�M�9��dr�w�����}��-򺹽�s���{`���V�7ּ:�l~J%:�C�4��bkdf���ݜ.���s�u6LH
��`���[�J�/�<J��Q�ĝt���ts�{��t'$�tF�ӛ'/ɢ�v����~")�:���� ��j�)@YʵoC-������~]硍�!���~k�	-��\��yBi�� �i��N�k�d�@�d�����Zݑ�0�4�Hb�zOt�͕GY(c�e�SML�I����K[���{m|�ۀ(n+F�`�Ԅ��H=�*���b��3�
ܧ{����֧WA���e.�I�ra��p_��i�s=���"Ƙ��&�N���`� ��.���n\��ӹp�kQ���e3R��~�8�df���mo�Yi��YC���垐#e,/o~s`�� ��+f]������	�h�?����!��\S�����<�y�^�=�n�ӑUo4k��D�)���S܎�Ro��oH/�7��~�������[��W��u`�R��~f���k40�ţ&���I��j/���ANB�٘��R�e�~	m5��^���:���r��0xx�^�-DS��	�ۥ�%i]�y����9������Gz|��RX�&������i'Q�׾�Y]g�V9�H\�6ZB:�^���֛J������t��ц3��ym��/���,0���fG�����J[�j�����1��Fg�l�=���)U-dQ3�A� ^K�#�� =�mU4_Q���Q*Q}o�kc�,Q,���R�}y&T���|�Y��G?)�n�j���%c�mW�}�����Y�?�'����L前Oe�G�"6�a����H{|���^]z�I���XK�v��9�f�t�Y�o ]��_D��������\����9�F�U0!�`2���V��_�������.3��Ҡ��C���G�^����ځ������F��+)��Y�<0 �,�5�W#x�з1
R�i3��/��W-N@NB���(m"ngH��rn5����tτN�.vƶ����s^0�7�W�d�Z���x��I�[�@�"�1�qm#�d-b�az~��=I&$6����1�{�'�s�dx|����T7|!~���T���{��}�dK�J���c�� q"������cd�[�!]57jt蓠�n(X]�ˉ��ل��t�������U$7YH����*(~(�Y�,���a�8�>��މB\X|�:F���K��zbQ���_s%5� �ԁ�|�2��Z�#e�O�j�D3�9'�j�[�|`�Vy�]����ϔ_��5�"�IVob��`'��&b�|�eE�^Ԯ�瘝D㼄n�s�/|L������z������� ��a��
�4KIa��3�0��q���9���m�:�6��~��K	}��ʒ���{#X	+;��R�@h�ϓɂ�{���o��2˗s<��t��_023��O�৞�9���(�ҜSP	 �G)Vq��	HE�ޔ �����{��6�Y������{�d��y��g�缌�򯙭 ��5K.�#L�.
Wd��D��XZçf�]���̕��Bpy]%�YQ�"Kg��b.���L�u�nΎ-]!SU](��!5�i�\��+�/��Z��FN�ʌ�`��n©�|�3'V@��y��m�G����밆螀�f�����Ƣ��5 %K����)U`ԋ��2QԢ��PTk��Fa-����f�I�=���#P5�O�"�ܘ�?��Z��j����Dtn�d�!gv�$����� �F�AC���.-��6o- sM�*���\ݚ�X�l�c�����)+�f�F���)b"����>�e����K���v��H"`kC�����57~���&�r�B�Y-H��0�Oί��l(º�?:I�$��V�[D�iL��]�zK_��m~`�T9�%VW�/|�XNx0,%�Jb����^��Wd	ء��f��m;����?�"��|ZU��R���'����\>bk�uQ ���)+R�"�:��]���?�@���.
�]�L�$�X���[/�����FK'�pn�����I4\�N�k��9W.��K����`�j�2N�̩��-�Rւl����N�I-为�ǁ����̸����V� L�ꀔJ^t58�D,;�9HY}b�R��9�=[c������N�so�ZC�&��-@w��,QC$f4a�;��&A�m%!��nW�L�m�Y��~�<3}`k$����L��S�}��|gS6�����K�R@Z�D]<<�\H�y׮]v0_�m�U�P� `R�BƄQ���?��'1jm���#2n�@����@�_��<�=����!�����"�/�u�$&x����SV�,J�=��
*j�;mF����BL$«�;�J"v�n���S�����1�h�1��r{��0��AII��-�,���Yz=/��W�-�,��;,�f�*�Ԧp����[�c\��Ȝ ٩b�T"� N��8��p����!�s���~iC"����f���&%��m����R�O�_�5~��_,%o~3��Et��6s&�mY
�L�#bn��ρ�O+]��Z�8�)���};��6���f�)��H���/x#��;9:8Ǟ2���E�I�����ր��?��%�E�?�[��>P{��/��W�R��,��'�F���zg�����5��~��$E�#;��9��΋��Mw@x'v�������ѳ�u�R�~s훫hG��U�ag7�x�c	�:b�]�i�_��}'2�\���P�`��O������.]E�XW��wߡ����HE`�!�ѱXvw{��~���k��w@
�,U� ����_��$f�ӆ_&&���ݠ�A/���M�����"�rY���[�R�	�6z0�{b��,��"I�Q�"�7�ՈҘ�_	Ŧ�/E@����O��5 '�����U
��c��k�Șk�����$��W@H�m!��qN8��ߐ�km_N�r�(� ���5�C4|ڔT9X�h�5o��{�C����ah�p�F�F�L�?w�����	����ŵ�C��d:��	,܆��+_�nm��깱EsWen�a#2{�o�.#sb��%V;Y��B�:?)p���{݆?T�/~�:ǋ9��;^3q߶2j�ۤ��G��XA=��y2�p�E$3���ύk��|W?�����gYP��;� �%P���G힢�6�_���+�&K�%�����5l�Q����{�E+/���9l���.�\��̂a��1<�6;פ������PN���+'�YPW�Ɵ��Qd]�=��W�A��^K���"2`uI �J�A>�p�JW�%����c��̍�W�#�nJ:ǶY@�l���>���*Zl���� k�w��2�n�/p^�x�Ri{�5}��0xx�F�`�N�
��c�����5"�F�ɐ���P��^�>�-����Iλ
H=Ǌ�7D�� n��:��ZlP3I:18���m�V�ѱ�X�I�o��W�	{�1x��nO�4ex�_�Z�����2D�@� /��h�2er~�@[ 2���e�J&���B tc��	+���uz�P�-]6��;tx�ى�SGP���k��Wt�sｺ��>�ނ�g�{8Pk��+5�y�jS�̋e�v�tb@�W<��Nh�<4]�L��
7H�+Y�AN ��,�i��+�t�4�1�Uv(���u��Oy��{��LXk�4L����d�>�%��*��P�z�b`��1_������u�_�y��������K$�����n��A%��<��r��tJ��L}�OH	�~1>`�>�	�+2Y�131zs�\bzN@��cL?�a�b������3�*WU7�8�*�o's�A5V3�>�s���q��?����M'�V���a�|m�gP4��K�~h�a2���>`?^@��
�B��tG��?�"�d�v�_l�;9�MO���N�ى�)������Ȱ9 {x������,zk|(��u�b��/�7��4d6�aܻZ(����<~lML8'!�C��y���nY��$�B�Ha�V�����^j��`n��&�3�s�}ß<��g��<��ˈ�	j�X�*}�"�
��@"��a��f���Q�/-�uqX���z��D`����kxACI,�����F8q(z̝x,�2(T$J�i=h6
ڜ�kuZ�ֆ)�85_7닢�֨����94��L4���
kQ��
����(Ӳ'/;ޛR6����E ��	S�:���;U��uA6^{$qn3Lt�� G��8���g��+�k+����W�w������܃�� �Y�IHQ/7�G�7�؏8�	YU�@�ߕ؋d9�g}�5�:3*ք;R[�D�u���꿜."]�����KA'����ϨX���ª52���%��Y3����4h<B�' hڸ'�3-]&�lA�u��X����z��<���%�TU�W��:n:�H����ǔ׬υ.*����'}��9H=��#�qĘ�#233�y��[���������o���5�x���
�nBc�n3��I�����׊�h���hS�c�W��-�a ����'W~ͦ1n8�%3}��S
�G�t�K}%>�^`3�B����&-��X�%� |���c�G,G���h�~�<R�Q��M�\Q��K^?o�K~*���N�Y�Փ�����2�9�?�3`��c�iG��_|q���e�A7�7����5��t������k�>߿�}+���G�=cd�qf�ɕ�~~�r0���b�	������t��#OZ��X8��{۵;{�sZ����yET\t~����*�ZX=.�~B�KiW��Dg\��/�� *$���I�1�aT�(�Eo��G�3�X���F��ײEU�3�o�um�o���X1Z�~}<x�F����7��c�5З;L��^���0گ��E�~����C�z�E�{*����[K5�uE	
�co88��'�p�rq��KF+SY����?I��w�~1�V 8�v	���åaF�E�7Kf���]���{(ģx�ڎ�����x&пbG����XY뢢J�S�4i���ג�tǱT�Vj�h�^��BU��L�~@�Z�or|�y��@�z IAܒ�x���>��y!K��1�clF��am$O�ۮ�u�.Q!�U�l���F��R��kh��� !�t���r!���4�
���^$P�ds��P�u;�9��_�pA��>)���~b_��C�@o�O��P�[�Eo�VhK���<�5������_��G���nɤ��{��̡Rz�u��f0�8�RD�S 5{�:53{&���m�2�F�{���,��i��-t*v.ǯ�
E�Tu�Uk��(�4��a�I�R���~�P��|��=z��_��FV�5P`$��+4~���1��k/���u(�@�Ϊ�Hv����Q��Vl�A�l�}��K� ����@��|�y��]\Ƒ����B2��+M0!H%��+��\����\��tX�K�t������?5BVyX�f|��$��(s�2e���o�����C8E����ⷌ�L}`'1g ����ԁ�Y-��i���BK�r0�;FX]���_�Z"�ɗ��X�Uc�)7-`�K�����ֳ�߲7����q�P9�N�4�b�2�k���ױ��������Q�y���A�����Ѹ���Xjd@�R�C�q��jݢ`T$��fe�s�G��4u�o��(����´<��aW+��"@�p�`)����f�	c d5�r]Έ���o�:�R�`�x�U_:擾t�?�RG���%h7X�E�Y���<A��V�;Y��KVZ֧x��3u�+���:�lIQ��3�|�G��
�=��&J��Ӯ-x:��^wx��݂���C�C��)��Kt5V����Ez��n�*ǯ���"��M�M�W���<be����-�i���qK�V��y�2O«���u���6�r*��Ҽ�\����ڱ+�nG�c���.9O�B���y��!�Н��k��q|�
�`�:�	uW�2����6Vt+��~f���p]0Z�%�M�ۑ{.ʌb�%�?֧��
2{�,�+ �~7��Vl_$v�֘;���ҙm-��7�ƈя|�K�}!�^˫�B��@׆0�b[x��t�[`��4FOx��/� �}��=�B�5C,o1�{�rӵ�3#~#�1�?���Q7��AĮ�X$�T�m��Z�`"A����e�S�f����2H�L�ÝS��H��G�N��	�c�e[���Zs����O)�L����#CW��[�v���b�T[u@����, @����RŘs4�/������Z�z�	Z�d�yk_?-l���z��&�o��U��f��Y��	̡��T�*/��G�f���+�0�/3�y���:����AxX�?U�X�9�N�	$�֤��h \�2U�Z�I�eA��+B�TG[�"i�* I�����H���.j�Q��H���]\Jz01����}���N$&����z�]4j����w�W?�! ���W�+��N�,����\������RD�&])��/D�F�����j�a�ZO���枈2�E�asMt+?� k���ji����T�x8��@kK��S�?G�a8��7c��Lc�����\��Ȕ�
,h��@uF9�e+�+'�d舖�u����V��nS�D��[t[�5MIԭ�z��Y@WZ�$a���I�0��:���{n7�,��5* y:�"]����8�oRPpw���`w*{๡���e:Ѥ=��������Qy�&f	��Z1�E�H��?]BS�:2�� �"��t�+M���0^���p̥�Ųb&���0�M��'��܃̅V�Tt6��0B_��ΐ᳉J�����T�Q�b�
Ѿ?��6M!0���2��tb��(�nE�c?�m����֔D`�[��^�l�z���攴d�0�c��!jf���ǽ�32�WKO؁�@C�2pڬ6�BX�и�7?7���N]-J�\�řg.��E��^}T0�@3=�B���s��kV�gXf�W�N��O����n���p��WTI&;2���ޜ�I;:�;����UnD�C;K�p�f�Vzm�r��K�ӟ��}c��O��*��dJ����)lLj��c�b��k��㮂Y�R-۱&V�ݑ�bR�'����$0������7+�1��`����bǀ�4E���v����G|�P�ܯ�9M��)�c�Ą����Abx�=�fD�7� ���gƂ�xz�J�݉��r�*�:;;��=�ǱWa9�@`�W�='�=f4d>�\{�\����1��(�:먪�ƍ+u	tD��tg��"#�B�w3*fB`D���-��O+���=��7���~���v�77f[�u |�/�%~؇�w���y�X$1��g�#�"�
��G�&���S���O� �hڊ((Q���T&!+��Й]�Z�ڙcDf ��8�hJ���ݛb5zh�hmZ��[�[g�߸�E���P��!Q]1�5�V�~���*��ۺ`��P��u�*[�+
����;i�6�sЀ��#4.�AB�+�l��Y�z��}��,`�~�I
J2�W�|�)�>5W7гsaʖh}h�%m��%tư�/½���01ȁ`~g�(岦y��������0ϱ�8��ZO�7b�G�L C>���3��N ��6��"������>B�@;x�=p���ş�tb�ɪ�yye�����*ȧ���\�35��?2ުfW�D��4�CFz��vt���^�����2��"T�5��
˂�8�"�j`s��v��7L5)��5�<�e���r5�k��������r�1+g��_���5�V��+�"��ӆ&�t���uK��Q�>
��y�������9���I��D�*@ǅ�0�=��*(�U(�{�F(ݵ��ˌH�=����hgqN���(s==���������4��\XZ���;)��|^z�5��ۗ�`/�K/��E���*ZW'�C\Dw�h@{`�es���A�/��3�y �Ź2�t��[���5>\�"�q����ٹ(��G�CY�A�4X�@�
���7�H�&���E�H~$��B�̵U�k>)�oO݅�����:�7��o�Ű�����}��ol}��ZJ���V��b�J�G�p.��F�Ӝ4�3�C���gy�
����!l�KQ6�-#7 �,W=�����A���췸�0��Y ��
K��F,���՟�������:Y�ΊUeja������=��Z��k��� �9�2x3��Y��j���2�&�xj�����W09�L�M'�r�jpC�����I`j�X(bN8��v�R��5�л����ҿ����w���JA����1�x���(H/RҞ���Ex1��7�G �*�Ot,��H���Y\�Ӊ!0�e��{���ļ����O�2s�d�%^ΪcD5��{��&�xu�E���k���lJV������}�"�
����E�#
͠�z<u �ʯ���Ѧ�����<+��!�X+���B��Y�
۔���	�Ko��(Q7x;,2��T0��c��/\���A�2�)�,��X0�A���/  S�f�*�������M]�������u�.��.Q����]��q��1��:�T��dʆ̀� �@�!a�ہP���w��Y�ۻ�g|�U vI<�W�lV�s��׀3�p�b�\IMך؟k7�>��f�B�T�'���j�7L�<ˠm@$�h�������c�#�g��m�Z��N�o��}�%���y���xa8���r��]m�.��M$ˈ��/�`�(���	�eKש�ϕ4@��\���8��F��:��"���u�����F��%�ei��ޗ��sR����a.��s��a]U��+.P@X���&���!�C��jB^`����I�d-�P
��O#V��,�t��w|�Q>�=.]�S�ص��%��Ӭ��v�q�������`r�M��)���<.�hlN/�#{`�JG-�A)9Ī1%��]��І(	:I�˰�Bvd�0�0��;�κN	��0-�M��3O�����@�����$��:����-�� P����P��K��h���^K:�A
�C�@1:�R*�fR?��v=�z�:���6�q9�_��͵Ⱦ��(�^��.U�d���� �im�!&�ĭG���\��OXA��S����9�o��a{|�j�g-�ݴ�Į	���Wg�#����e�w��vG끅�1_���j�X��V}�R�^|"Ѕ�����F��Kc��˗C}�0����G����ʌ�b�U�0>�j�\���NO�˜���c6-�:�6#�)��I��xr/S�n�|��V�=�o�����?��|=R1ٙ���n�U8���%T�eK�ʆ�;�~s�~��Ɯ�U������Q�JF��⩣��W)_1=�j'4�
\�����@#efgU�@��b�5b 	�+']?��~,�i���X >:�k�ʫφ)K�43�؝kg1�R��&�������<�SW�;�@,s�	ۭ�]�ELW��]|�ؗֈ�������O�TL(ሻn+�"����v�~z?��̛=	rF�R��K8pC��G�N�aQ��Q�d:���H4��SK��ۧ��g���F���	���0�������.�[TW�ɻ��ɷ}ձJ��Ho142�4��ѻI ��W��->��Q~��J2�F�Kx�Y�ƚ�R9S27��}��v��L/]�࢞K?y�rB܉���Q�3��p:{��% /��fϤs��W�>|Iޒ��.���Xu��~�DfK$ 0���X�c��qP5�[��ދc`N�p��bB�C���*fּa����dw�)L_��&�m|q!�}�¤T��\A���Nf���dr�;e�d��7�4MT.��Yl��]�^0W)aW���;�=w�Z����()�XJ׍����+~u��N
�9�MkaǹM�Ǿ������ڞy{b{b�r�&l��|���h@ޗ���������0����
�O|���XR��؊Џ��������,6��ƾ4J|�ޑM1�fU�ǚ��b�FYۧp��_�&��ˬE!�B��/������mǩ��u  ��غ��|�T��q)s�z7��\i^'��U_C�ٔ��7m���I}�=��a1VB�1��j_p]܀Q���{��$�/DF�G�l�k�.��Ȗʦ�t��R��\\59�/3���'����R�b��}kDrC(�b�H�i���U/+��Q�:,$��+��?��m�(�of�����_،޷�~C[��^��ֽ�m�Ro0I���G�L���Ru�����G�ؙ��tg	��&��,��%�z�;�.��tE9�	}(����t��P��� G}jjY�(�'��n��V|7�bۃ�|%��O�`��޾�-*�=Z�=2�ݠO��������������j�@'x�4����A�%�	�b�2���G������w_Y���Mw1���ݷ$)�@��  ��ЏM�76����K�\q1p���Ll<b���Te��R |sp�_'�=pg��9����`�,������~���� �)�'a��>�bC�!f�A��܊a]�8�=�7 �z/��L��A�B=b?��琱�'�
"��G�!~��)�j��)k�}���y3Ԫ�0�%�ǞS!��wX[8�a\G֋ǀA|A�*r�����}F+m�Е�Gr{r�
S�MV|��G"`%�J-)fo�bu�����][f�8>�_DG$ �r�3eZ���2l��G��aD*�f�Y��Y�"&���eH�?7�ss��h��J��v5�b�Z�O�F�:Z:o\�8p�ފ�����Ksĕw|�,����"�&� W�vo����)�)#��Q
����ш����sXU�ʖM IQ!¯R�Z7t��������Q!��P2Z��~���]=��ÀY��{�`��b��K[��R<���I����&MQ^_��j���0��kQ�RK�1>���
S�~*�� �[���0�=
ZƼLR����9*PY;�~����E`���<�����qV؃Y�~�_ n��z�>P�5
���Kѥ`1��-̸���|��
���#��OU$D7�L�+�d��9��N�^�B���d�i)l�d��p�����O���]���3�t��ġ���(io�N�E�#2R
�)uD[b�I�m'0	��]O1��u����~S}1>;���wR%X�`�C1�A�Z�\���vHFD���?y�)�J�!dkt�5nt󭋨�����w����0U���LqZ����df7Mw�?Ǖ�����^��ӫ0�Ӝ�����W$.G�v�4Z���A%y_�_��;h�.G��c�M�/����hJN�4�p����)��;{ h�s�@��K�����h��A=�J�|#?zib�رl��.�������~��6oƮ��r��ߣ�OD�0+fg����K`s���L1X���<Ĵlk�N��z�)ۢ�:8J��}��K�v +�;JXh&)3=��4�̂D�C�*�ЬCpgaK(�U()lW�X��hq�+:AN`-�]v����Ǯ�Iht�Q!��:ox5�/���,��ϴ�X�Z��Y� �_x�e�%w��O����oa�I+�e���G{�̶�:� #sR�>o��N���/����߹��F`4	ˉ�y���k���}��M��ypX�[<t�B�^�����0�!���p�B�ۤϋ8���ߍ���8q$J�3��DU��5��A��=u��ya;Һ�>�<�xإ���~v���ۖ<ԉN��6�ҏ�.F#
@]�d.�PB����p@uh��<���܏`k�2���SvV�� ��2�����&I	�=ϴ��t9Fݮj}K��D�|u$a�m����$λ�K�"�A����10���5���W��;{Q�LΒw6�Ѝ�h��u�Tc6���$�0�$�K8N�2��}�d�}��w�i�'S�^❩I�Ym���0d�)��Y�E y0�<ZjY��{;���$M��xX���{nU���<��@��4B�i�{��ߤVX�7]�4�_�:P����Ki��B�k���an�=�������8�K��\�1Pt��Ž��T��9��#��I�����K\�k��ʩfq��Q�K%��vv��q/���� � �@��v��t��ZE��d,@�0wZ�����<ge7��+\�F7|�E�3}y�����T�,���jn��٣�0���z�ɪ�~��dyW�k���m���(>�R:y��&8m�,Fq�&���_��@���U1��J�_�?�����	�9E�Ϯ����)��׳��`'�i/E�@n#�47s�Y;��.���R*�f��CXs���f$瓷 c�@M��YbS����7;�:���K`!a		J�ak��$T�u�>�ĉ0�d�޷r�����K��=��.���oL�>��@�������AU�	p�T��;��I,����G���x�.���%;1�5S�� -$:H�?�s'V������&&f�=k�$
��ֻL�4�:���*ҡ�F ��<���lS�sM���1���3Ӗ�l�����S';�_>������J���_(]�:ꜧ@W� 31c�q��v�M�Rn�]�ƚd��d<p|���SB�X�sL�<>la��-�p�;�b�� I��g9L�~��Ί%׹-��@�N�h�M�l��Q\g{�H�ߞgJ��5ƞ�1\��Ii�T;@�⌸���A��-e�Q�����_�&�Y%�N�˿^�,��?/>26�=w\�����1T��O��JV�����1��,���)��:T�����O	���</�l3��+���a`��`f�no<f� �	[`)P�n�iȻ�0��4K}��� �l���������0�n�m*$\����SJ��o�o	7-��\�J�.�+�6� G�-_h��Y9^��5G�Si��O$�*���u33�?X�@̧J,+~�{>P%J*l��H��K��(Nw���8��An~�y�|ՠ�dIr�XȦ�1�������4�~{V�~�QɕN�.ě��2��b�����l�.;��(�P6��%l��� t��Ϻ�jr#��wͧp@�� ��jDf�����t=�ٜ,�m��u�L��o�C�6�u�)�C"N�d\�i������JV�F:< DF��DZM6�^�9��}���Xb�m�ֽ*#��3t�a��������>:z�}�� -v,�x1��!8��3_��cǯ��.e��W�#�J�n�DxC�+��Jʍ��,����i��$eYU<u"^��ɳ�X�Ǒ��؏�r"/���D	
�vԈ�X7�Y.H4k�r���(`V��
�ʐԴ�	R��WSv-�S��{�z��/!��۫[�[2�e����X۶�/���(�Z\�z�繠h ��L��4��6N�-��D��J����;C���hټ�_�Y��|;\��
�������0ٲ�=���� �D�8��X��8C���8���7M�@�y�6Vb����4�Y���߈,WO.�'Ӫ_�eUb{3����[:�ҕ�y��.��oL[Þ�P�q�f�oݽZu���r#���ɞ�9)�!�v/D-�	�������yD tpf=�^����t��xC)�dO�Β�x�f㱆��v�e��e���	�~
���A��#/-�SB�Ɍ�^�x�{	�C$Gg"�_�t qR�O5����Q�)�Ug8��=<I��b|6h���b�Ԩ����	������'�n�r�ݶX���r�ۅ�%'�w�J
��9�H���1*2�/��''��ktDy�Z�~7��86��d/�^�!�P���Sǰ39v���s�H�	�� $�������C*����}G;���Zu��=��S��4�U?�̤����$vce�5�ȒG���L�����<�5?3t��A����TR<�숌T�g(�?�����;z�5���7�� &���a�-؆�pz�q=F�� o�=��s��aA�o
;��f#"��0�qd,+��Kw�5���G�1T���1$�~E�B̭�6M�
k�|������-�Q�E7)V���}���T�����Tٱ��&d���
S�V���G��U��
-�{�gz[%�&��)K�su�O�j>���<����	���$������$�����Vz ��<��Ǌ��>��}��쑅*։Jv�bc�~�4���^����g�2-ea�*�vzu�M��% �>\��V���
�Q��܇P:�lh^�=���_��*0�h�*�[�c�|�E0�#0}u��D_Q���Ye�"4���@��{�L@4d���*Aa�q�3>&��>άI�����2qr��=9�!�����g��������W`z���n��W���ܳ�T����PWfEtAP�2��y�ͺ`��F&�T-�*�?���������{iN*�w��⊲tÐ:���/�cNe��EB��N�,��K��8�cg�/U�ϣ��uk�4��%`e7|"ޭ��}����u5:��w/�>=�.P:WLN�N��`�>sJ�dD�Vi=XDvS(�Z]��|'9��\�,P�� ����Q&�л�(�5,������"tM��� ��Q�y�/v4��sy��lF��O��Ud �د峀5��@J��ڥ���8es@=_��ؘ	A@	���9�-!�U�U��DA1�o6S-?�h�M0(��n�-1��j3t�ތ�\���V������Ɔ������3��u\`	��#�������E����foI	,���M�/�m̟�#M0�%o�<�l}z*nR�њ2�\z�3m�ue�dX��6�K�E����| SaI���]F���3�Я N'y����9�
����Ǿ�p~�R�;��>953�;�I���dE�x_�P� �]N�T�������ʂ�M�X_�k�}���C����_�{0�h{6�R�%������4�(ᕜ��{�� ���}��%bh�$���ұg�_d����Gz}�xo�sq����(�{��f
�^�Ζm4(�I����������A�QI_}>�"��E�s�Y-�ǠI@6�[kwʻfaJ6����=�X%20!u�e�� ߑL��3I��5�D�-�X~:�n����Z*VT����j�@/�{0
Q ��3M�m~X�3�z��͍�E�_�� I6|������)�n��Č-B(��4����]���b��?��_����I����J�2쟲��}2n�A�>51&-��CP��p�����a`�K ��� n��"��?�`W�������x��_�G7e�	����<���x��n��)�OZ�ᶔ:��/1C���Z����*�k���/؈�d޺��R���X�[ʺ�Mh���%Α3�e*+Ǉ�<I>�0nz���:��[�0#I�[��?��7W��Z��(�w��P���b�tب���&���s*Dx0{�n|@�[U�V�Z�R���gvN�$%� ҙ�1$M��8���2]y셏K.qp8Z]�gMpPݵ^���89E�K�ZQ�h0�_)�:uJi�|�s�*ƈTc^��"�,}(K�^h#���ޭ�p+3my�I
��}�ZG�S���9?�Cx_��xE?��(y%�EoHe�R�P�BKA�o�yοO$�}�͝Buc8JK ���!ľ.Ҕ��֖	Ep߾r�%����[U�;A�yH�Z�{7�_󋾾��+��=��^���.^{1����b��{����R��tcH*��R�/Ѵ�'���|���opJ����3Gp�r�+�E&������� ���/�j`T�9��C�26<��Y=-gL�i����!�b�����C��DTɧ�`�8WW!%�P������,�/�X����$��%*c�m��W ����>=��1J��ij��y݌O��%���bTϚO�ô������Zأ����it���tq�������i�GhK�TU<sa�`~,�}��8����m�o���ā����\-��L�6$=W����)�0��V`��&��8��&�(�	�Ɲ+�����"���)��B�ϡ� �4�{�A�',u֔�qc�@զ@��:3��5�k�f�,��1�L_�5�DQ�ᪧ�f96� �w����uΈ�u\�'��ߴ�<�Q]܇ZX!ʤv~����Q����A^�aa�U;�MH=`��0ӻ�m�AI�&��T�AZͅЛZ6<s.U���=�1L�aaVZ����Lz�����9�B��H� mN�rnά�F.�sI��<E�� �Z����5��gR�oL������#B/⶯GT7b,l$c\?j����N3ov�y<���K�۱�ۛ��TX������n�:���ר"9)���t7�o��=�u��z��}4�_P{j�N,W�Sg�LL?!�C:� � IW�v�o��t��e^L���a��e���C����hp��SN%��PP��u͓�죄T�%�䯐~���p�`V�G�CJ������=ς�@�j�	����M9?~_�#k�G�>���H�w -H�G?O�[����?%�Y�笣��?k�5�~�d��]F�Т/ӽU/+������jk^�n	H[@ߛ��7����@ro�9S5ecJR �[�Vx��j����e���\�2��lTA��ߑ��S���p���>��cU��kw����P����eXf��6{	G�/Wd�SF���|�%�;'C��S�R�f6����x��,JA�~*^4�EVr�v�h�����������Q)�RjM5'���\�U�z�� ��$��iq`
f3w׈�m�n�]W`��,��.���~�(�?0�b�ы��Ø�l�
z,Sht.{�$�����f�	���|9��.5���F�ҖL�p«S-�����q���w|S齎���w�exL��J�Q`�� �[��l1@�pTr�"Z)�'{��_�X9��o���B>�q1At�?�,EݧF�%f�K{x����o�M�G��ӎDK���a<N�y�;����1<�^�3U���.�%9��=h��Ӥ�Z�]֩���R|�Y]������I!�`���"�E�-��Uw�=�5��F�	G,WD'[R�,A���|�ފd�f6][�^q������'����Y)-��ڂO�}�6���0����lG��n�b����6q+����*:j��+�CT�A�K�&G�hJn\�|k�%O��`k&��Y��]�/Sʺ2y��T/3!�L�����C�踩p@ν���J%���bpQ0�'W���[��,��A�H`�>c����p�9r(��{lM���"K-�6��+E�̙ݠ'q�R�ހ��wӲxV�0�&V�a�YŨzw5�g�8m~���On\����!bW+�:}q��]��흓Þ���?lI�l�|�PuG{�����h��7�,2���]dȾˍ�@�L��o�M��[�o�R�;���:�J�����}�2���3�Ȃ��]�v-�_��Hx�I?�ᾊ���Td[_�l7���H�1��d�nO�Px�j�ףqZ�����t�e����($"��-�>������Oqf,쿓�Ŀ����jَ�[�֬�͏	�Q��v]�⎼ne���M���M;�RQv$R�e�Ä�����Լ�2#�,�����M�cߵK�0���ͣ(���N�d�8%�Ԍ����.�$~M�Up��SHz��`7f��G�����9>��������f��-Ew^���ĉ7����.TT�_�Ҍa?�!ә�a"���9уs�G�m���yé�e�ձb��r/H���+��W��I'6$�0��i�_�9I�n'~�z�;}�է����~��^˻v������e�iN����c�����Bd*�T?���OA��aɡ�_�T&�ML��婸G���sv����r���̶��E��QD�Q�t��d��Z�z�^!,�1���e9Ξ��֯6ܧ ��~=@��Ph�#��3Q��F��N]�?i�<J��c;��ߩJ�@D4k=
`�|���F�(���|}��޼�^��<�m?���Q{����H�{Xx���I�	k��װ[W?�NUx�f�ȹ�g�ȃ��|t��|�yA�G����;���.�����L]g@SK�zp�WT�#]����H�%@�*R�HU��T��� ���*]BQB�Є�B�s�����_����g�yf��l�5�ʟU�����&IN�Ck�����~r�}EkĎ?/n�SU�����荗����X��7���[w"p���JzL;�^�"���ފ�j��`I�;��z���R����(S[Hș�Wӱv�xq��*K:k���#�1/ialU?���3����	���C\�d�򡶹>��\I5Ë:��Zx�bП�x-�#C�τE��:�E;A��A��!*��Rj��2��H%��/���,���%M�f&�:g?�,�B�F�CD�1Ĳ��oNm���h=Gm��f�Xv���S�0�Deݭ��P5��.�ZC���0�5���ӟW�pդ��E`���\�`�+����[�_L�/W��s4�u�p%�tj���ꃡ��<�aL�L�8m�����������<���Ǔ��,�¡չ=К>�(շ$�����F'�<CG����`ӛ��_�����|��%���ak0�X&6|�a��ҀxQc�𔲋�/d\�j�S�K#)h%�le��[-8��s;�^`%���9D���w�hzuJvP��UX���vJ���{j����w�{��?���,���w?�ΆPY���w�[ pgW/�F�à�&|��c�h��{�J�*N2q�JR}p��OwkON�S�����|%�c�_9�5�ܘ��-�㿙7q�H�L�G:���'U1i�C�x<�Y�����i��n���w� ��V�z�Q0j�����9�����C���Y�z"4D1Kv�x�8�b:�;Ow"o=�ey�ѬL����2���������v�,��q5W0G"��,�c�,H~���Y�=c��^������Z��Y�ŽmG�[�IX*�y+����N�k�2E�2C	R���b�������"BjI��+P��O��v�d��F[�����/�Q�N6�BO(���p�j�q����TNI�De{|��]�q�	����_dw��/����[��m����d.������d���W�G��
�� Ȼ�k��/��Rv��~�����p�1����PA��'O�Y���`�Ef��ӧ��^��3�^����ͲK�oM�@5��im%4�C��٫0��T?W!()	j,iF`:�dW��aQ/���k�S���R�����S�/�:Q��z�~��_ӘO��hN�B����w�臒/�3(��%�]���}������l�;S����6�#��OR�2���)Kfd$�[����Ǝ�M8��)Rᡄ?�*[L�$'�tL�-��d���$�oX  =��w��7���Y���jK��qP{�s��h�R�ehȍ�w�q 	ժ1ۅ���rL�.o:�դ)[*�P��QO%�`��O��HH �F�ͤe5�Q�p/���b3	���EHL�#n�{.��FD�do۹?�j�����<$2�CO���kE*�~�����Y��Crá���/M�k�gቢ��/:ܥ��82�I=q�ܨ�#���my��Q�~S�\2(��`:��p� �wH����UR��j�nOB�CO5��[K�\5}��6^�ýt��Gv2U�=��rM��mԺ��K��ˎ�rF_|��Jz��bה�,ڹI��ڷEY8s��˗]̤w>�b�@��r�H/j�iLY������&�r������l�ܝH1n�R�~;
״���KL�Qo]e�[TVx���Z�3�l�V�����2U�
��g����I���:�w�4ńN���;*��.1�>4��{�LLf�잦|��7�|8ו�*��X�qys����F<�n��@A�M�0g����p���j��c��֛�N��}�'
y!r��ñ�x�4a�RH���5�<���kQ�i��]a;�ұ�ר�zxv���G��\���0�J5�!��Gn1\[�{Wlne� �ֈ63力������:�j�A��,��nZ4��:B��!��~�s��E6��~���k9���q���)�uAuQ�Bߴ�w��s�}�'�'���1S\�����t�s×r���IGs�!?�o��n_Mk��l$<�YX#q��F,��V'�gT�O'3������홚S'��u�:�o[xڂ�֪�nb��+$3������G/��y_3�|a�[TS��^͕l�<m ګ�Ng݅�-��b��ܧ�aGX+B|�``��dm4��^p�.b�o��B��S5��B=��C�4�J~�_ۚ�",���th����]�$�v��c���n�P8d��?7���`��r	�R[�;E*f�M�F�R���e�M�����K�\j����/�����9 ��)h���r��T�����.$�4�nLn��¹�����*1��?����s��e��{eQ��S��l�����|����,!�:�{�~o!�J�e�Ulg�FV�>Io��0�W3��9Xp���ҽ�m����(�^&E]��-�*�{���4��nǔJ1S���
6����8΃�߇B|B��T~�@_D�a%o�������exa�����.D|�(�r��Q	�~���~�z��0������@�?T̀�t��i�.��x�2,)����q�6�~V��:�g�S�+�J`U����������B��I��Q�;/�wj	����*� ��̝�.�f�c���'����졧����K=��/���'~�͝:ع�͌������Oy��8�����H�!)|�{�uS���$�t;-�:����.�X?�=�,^Xmdˏ"�=���y���j<G���A0�<��d8����������#��MUbp� �irgP�Wv&���_�Ty{����Ub�a Csc�
�mK�F�"������lV�(���X?���f�e�j]#�c�}a�k`3� S��%��T{7��z{������j;)��&�[u@�ؘA���܏ˑu5R���<-}� l߻��(^�tW6�&,�*����{��R�ù��g�����&�k�Hy%y@v9S׹�+�X��]!�rݗ"�Dn�ٔ,尞��.�T�v�j���9f� R-{�폿F����"���h�rs��5��{�$��6{��🙏�<>z���i���&7g������z���$�2z�V�a\�i�_"����^�D��!�=p$#Ƽ#�Y�5�;�ʥu�DR���3��\y�Nuk"��J���ߔ�b]��	������� U�:�ͺ� �OR�FKLב�2�{(S��)���,�6��4�Epq2Q�����ґM��&yl]� �9�F�a�ȥ���8�d����>�:���=�9�5��R�nkF&�i竷?b(�4n�IM����FU&��'��Jz��E�{ y�6���7�L~��[d�0'��tXVb`���(���Q8/�����K�Y���b��6J��6a�C�в.aN0l(����0��F$%��)w��4A�C!"
��g�ٱQ]�j��O:ʮR��SZ���(��j��<�����M9�]m94�!rlA��U����M�YC�Ő�N�ڊR�d)�j����BOdꩄ�����y�wI�/�A?0�暆x��j)�~�F��K��r׍���w.,�P<靬��������� ���l}����#�2�u�x��;t�T�@پS�q�q����A�܁Ef��|���l�׀Ph.��h�\��F�g�۫.�r&a������-r�\X����t�0M�iD�v�@�*�|y	��]�MO8?^�H辐�6&(.\OpM��e&���0}��L9n�F�j�����Zy��(?��!iy�g*��u��]��A�H!�{�d�};L����'��_��6�|�z�#�R#�C'�ö��F��&"�+Q�&^��@�I��1P>��N���2n`0�Nh�q�8�A[Š��9,*rf#��3,C� Ȟ]UW<~������j��hZ�����)�)Z��+ǜ�����閕�����
�J- ����m�a]&&�*)��^��g.�5�S�(�uR��y=�3����Wz��Op��LR*]
�F4X	8�᡽[�Cjʳ.#�A����Jg�f�|8���m���`$���\����Մ��/@(��髊��B{�81��,eg:ږ��^ؓk�����)>½qw_qcLy�7ִ�����*�F+�_�Nz$���%P�bܡ�mQh�{�QH1L�Kr��G.;JVPP�ӻ7�d?nw����)���G쎢��:��8q[ա��@���##t�~((5��Zb���g�=�]
���:!T.ܨf|~����["e����L3_��s�=�$=E7&��m��w������4]�wvDu�Q�Qo����(wJg�a�'MS��rW|h��?���ri>!���#���U��j�k�.���x��ZW1`�9y�x?��Iʩ����yR��g���P� 
̋��5����/ov��+X�Fp���^��؀��=�T]נ����)��T��.0
v�����L�)�Jn_S�hn:S�(}���eV7�J�F�uj��;����kzG���nρ�����g#��{�pW���������("��S�n�O��r#��0�� mM��
����<g*\2�Cʪ��t���1̸RQt|p�DT�����9�.����l���2�m�{�4"C^^uN�j��� z-�mexlnC�,Ě�mM�	�2~%t@}�#T���1ԕ�� ��2%��v�>hD{��m���9����0})*���ٸEr�ۯ�_w���lqj��L`�2�#���7�����8�Zbo��!�"�lI�Q������p9�f���z�h�:�3T:^�%i���CL���V��I�f �����
 ?�V� ���ٯ��������"j�J�j�1`�+OU]�	���&��$���o� �>�r��ӫ��:T0����{�q�[!A����P�S��B_5��	�.\.x-�,��&�cQA�۩<ˏ�D�t�����x�}�;Y,��s��,�&y�_���2��`_���������0ec@����U���)��az��ś��DG����z�@?��n�ݬ� �*1c`����|���U=]����>�z$ʏ8D�O����1�L�Y��pTh�s�؞vL�z��2���Ӳ�,8������ah��z;���������rz���e�$ߧD?�z�qAXJU2�4�xSx����ԣZ[,v_�E<���A|�T �*m:^�p��B�+<�]NԵ$�E%����1fU�1!�8ꦵ RWQF�P@���['�z�{����L\�g�Pu��r�MExkOB����aJ�xi35˒�D��&%�Q>o��]����j��r�vmI���-{�tN��_i��.p�c�*IN�(v��=�K��4���{1�� ~� ���N�MNޱ��֡��,yv�o�%�<땘eQ�n��Aj���E%���:_�t[�|l������ش&�m=KrI]"�J2���v.����/B5�>�����D:�*�ѵ����cB�3��j��
-�md���F�w��SAv/�D��y`�X�BST����H{���y���G.�:z�r�Ʒ{�[q
�g<7�N8�r��V�����?_��=	��aJϺ*C_�k�J���2�O�	������N��w ������_V�ߌ3z��#Ǥ&��T{����[;�q��do��M��nRC�@���i�U���&����>k7�\pB�>���	?r#3͇'N��!�g8�S�2�+�;�h޵�M�.�1㹕z����% F���V���F��Kn��H�<�*�����.{K/jq;Jͤ�Zp��I�`�}��3�/�veZx��g�� ��XL(��	g�P}�/�?$u�KWn�x�neMyG�6���j7<��C��i�n�:TmE�y�
�"�����Y�DR~/����	쓜�7ZN���ݪ�u�_�A�+<m#	.W�*��[U���k�/#?����|E n�������P&8}ڴ���١^�T-��_�CC�'5�(�������8r.����p���0h=���"W?��九92j�Q	�`#8��j��:&4J�^]�Lv�ڮ"�^`2�}YnKy�`����j�����,3�f{�+���\�"2n�^(��}M���΢�}�ۀ��8��p����
�Qe`5m�������M�򑬲�	�K+�����%H��q�É�����,�X�K�7�lPsç�څY�
%K���K7�����r���k�5�|���������X�>s�V��m�&2i��Y�>f���j�[M�QS�����ޠ.H�ʻ��[ėԺ�c�D�2�[��F�MI�4[��G�ؤ�
e^k���'�H�)M�1h3��YL!�J~d��#���i�hu���l��GF$��|��]U�(�4h�2��ת�:����P]cW����9��3���N�QI�G�L�dW'����˛�C#���N�\v��O\�?9���_���¸FX���Ϭ%�]��g���eO�a���	YJC�Т8ز!@�Zʟ�,�HK�	>�nJ<��$������y�W�`M�HSf<���a#���gx��P�^$�~6�-(74��FI1y3Ћ�gc9������+]�-�0W0�F$wΠJ��� ����e�N���|Q��m�]�jS��$
���C����j�2����/9�G���i�z77�J3�|I��̘��KD�����*����#��d����1�c��M�6nfk��y:|�f�慽���{G���lYa¼�9����痍��e����A�nGnj���G�\YS
����r�˸���������z�|���PY��~L�,[�u�Ӎ��z��2)4���}�c�7���"#u��4(XD����W�gs��Ն��Y�渽_���T�1�(�,�M�u��n������9 #���,�����Z�3���FB���o��IĬ8�dx��e�]�ɗ�.����Ӹqw�:�j��DͷM�gHс!^rݠj��W*���RTf�G_.k�qs�P�rØ�5���W*��,�}߷��%~ ����;��u3�9yJ~^}�ߨP����1��*�%[�6d�q�ɼ88�}���l�@,p�qP��l�;L�C�Y6���������C�{9�����oR3)���v�������l�_Բ�z�6����>�Qg��;0�6*R��P$q�CTJ(�W�iŐ�>n	�#T�O�0}3ں����0�=������5:�y@�d�&P� �ƻT��)�R5䗖�r���X������U�Z�o�p�e-��z�ㄇ��J,�����N�Z$���a>�G>��?M+_a9��Ѥ��\ڼnĂ�-	�M���Ɨ�3��8��^,������v�R��f�/�W���C�F7��}Ɨ���Mi�
)�ZZC�}��(�C��eٵ*_��~�oOIs?�Q�k:��f�!��b��^�d�Y�x�AQd�2�\�	�K�1|�,<'&�IPG��{���c9�o�Nyp���pA6��國�rp}o�ދA��ܢ�-��z�;�d�*�� 8)�Ƃ\
I��[&��ܬ:3D�E�lne�i�ť�]5�18۵��L#?��6��f��t+ �E����*���"���b����?�e�!��3��v0������0���nￛ"U��X���6���l���E�h� �b��4�c�>q�R�#ұ�g��Mr�:,9K� W�(n%,P�U�ۭkO[6C��vEwx�����K�)�k�^��:�fB�D��[$hKM��m���L�d	���\��u�gX�(�Pi!�d�������T�3BnrM��4n0�n�.w�[e��c�G�긆_�Ҿ���I|�;w3��rQwb��ln��0_��@��Y�Qu�o�x����<3�����R2�aBh��X��ݖEn2���(�epdT0��(�.:�A�˲�_�}�4-��P�	[��"�R�@Y�=?ˇ���L����d��G�tϘ��B�kD�|�J�1)�]?�k���T(1�8r���͘�[_�姧Y�J��o�w��� )ȕkn����+��)Ϳ���+DV.2Ⱥ��od����I���G�o��MQ�oˢ��8��1�JJ@���==fQ�����+�\	�x��gW$}M�V�'+n��2 ��ضi_�?�j@��1;Q�e~�,�=�vX����Dc��+�!@�W�7́����]��GG�� o*�\�E��4 ^-�p��`�j��綛���g���Ik�kqN"!y*�۫������M�hXq3�������LU/y4ÂWsbb��3���""\�jo��T����<�?03�0�|�ċ޺L�q���ejw[�bej�0�f�|���mI�$s&���l-<x��Q����Q���f��\�ࢥ��^rrm�H����n�@�٣R0���U���I�?�S`Zn\/�vhls����xteed�3S�|ߺ�ұi��@,|1'\�2h�b����!n7�������O�P�ݫ�XZ�����Ր�Q�Uh��8 �[K�����WVG��ip��Y��ay˽
R�h�oX�� �Z�f��Hi�\,9� �"�Qt��9S �"�����BYt'c�ٴL"�DR<�J=�9z��P
]�/$mT��h�����w�7|=IN;�MXk�T�)ﺆ݃�f��.����7e�V���>�Z*A�l�=;ԩ�:|�=�����J�M^d��J��Zښ̴�s:=�5��p`���Ȱ�T�3�����%�O:�ԭ�o=2�o[�p��d�x�`�)]L�<G��	(R���v���)p];��4�4j)L�&ni�~I�5b��j�M�`����}���鞞^77�@-���Z��XN�u�Sƀ޵�=}�1�<��'�X��ĳ�~�D�1�-Z*C�$I^8��UT�^Z�?�eb�|�%�?}�4koi(h�K�pZ��ucHYz&�Z�ɮ�h
�"d[��=����'�@p��-���VA����ժ�����IC�����:6�g� ����v�*�i͚O�OK/�?@�Ȍ6s�jR�念\cֈ�si>�,m��ѓ�)5�����Y������Eù�=����{k��a�j(t�	���R��j��K6HWٴhZ�����9����}
�G>M�=Q�ӳ�q���y<�⡱�Yx��EFOq�N��	��n<�:��r��K>�Q=uܲ�(�Nr��I# �rD��R�i%���կ���UC��Eg<�
��@��H��"��Va�J���}᭐ІM�����<�&��2�H�ť-��n'��s��嗇�t��-�H�\:�1�(\7����ď�V�^|�%ZǑvN`�ʥ}��Y��Jwu`$�M��GH[�/5[hu�ʹ5��0P��m�� 0��t���e�ǐS휜�˸)\]��`˸�]Q�������/��h��i<b�'��vdAG���+��h�í���q���e�%��l^I?��H��r#N�+�`�w�W�TJ�T(�t ox�S|(��*���H	G�f<�蛉�ͣ@�6U�S�#��!�tX�q�B��S{E��mu�l��˧�&d��?V\���՜�_)�S>vr4=�'3���H�MԆ������j������z�M~��OSx�jy�֣�G��m��0��cy�XB��Ǹ^,>�l��I���E:y��rǙw�<����s��%�o�s<���ETiD^R�o/��Z��WF�7�	<�t{-2@��:�V��Ώ�5�["��a���6M�]����W;����}�rC��=��<���B����T�~뾢��+Ktg����³h�9����+$��\��!�2�S�w"�D��u�m�=�Ğ]��V�ĵ���cl�6t\2��A&+���< �[��f����6�@�����q3��q���!��߇��τ�.
B,���NdJx5�>�����s�9�i��C���v��l�0��3�۲rV�����!�l<x���隥�쐊6���=I�6��~Z�#�
OZ�'��2C˹���W$+���z:.ӮJ��!�>�W��𦸵ȟ��]�7;�r3v�9�f�ˬH��\�P�^��䰾�#�;�w��B���&n�������i=�q�V�}��"$Y͑O3�M��c;2<��\.�Q�3@J޻�:��m�.�:Bg���E��b����n�'���)�Ma}�Y_z+��:gW�~O	�����ًɿt� A�7ɘ͸:GH�L0�8�,�4���"�tzYr���V,\n���+ �D� -^J�4-�:�ݯj�*/̥��3��a��L���c8Mw�"�0����n0*��/�=3[��`����m�Q�@RL�����5���w�`jøn� ˓���t����t�뷘_Ѿ����ʼ�r��{���j+�٠��m�0g�2��|�w|xhP���FS��>�ҵ���i�["K yzP�&��q�=�����G?��yK�Y���)n����0C8����J��/{�� 'Ɍ:-\Y8�O ���N�B�
���sz����c3-�F���Ua\;oh���YeUO�f{�	&�O��ٶ��"��Sސ�ָ�{&�x�Ǜ�׽������9:-x&�;�V�k� ӓ���4QS4�rP�$�*ll(��IK��]?�R���ȓ��*�W�G=+�Wl6P]n[zl��J̔C]�=���*X{r��FjLaC�<�K��v�0�j�|4��|�K�����>�����m����J~�Di��f�!�P�q��3��5�T�
>��bJ
����W=�	��=q�8�7���6��K`��U�m�T�0�B��x�m���>V���@�CZ��2���f��+�)\˯n���|�f�_s����̳����@h`.�k�X����~j�/Q�5��&��c�������A?�4���e�|\���M߱�0�vN���2d$K\2#Xks}Jz�n(�$���d=p#=�I�i~.�yb#��v�w4��{`�3�tI"N*˒*5&��U�9��h�n��_�0	���� Pzu\�lWn/h�-�,����14�R^u�����q�h4��6mR{6�/ņa
�qkc���ר�r�(��y ��-%1˯4'];�4S��wJ���2K�l��@P���Az4f���H�)�  ��c��UP�c�%�V|fy�j��nn�^,n��bR����u�ྼ�*N�}4dEyU�_7�.��{O]�>݃�8��*>��Mw��?�J��kb�{�t9����� 5e�(i?(��:ވ���TmuB��Ƅ�����YՊ�6�_��tF��̯c��R,Ym9���{��O 6����t�	y\�ԧ!n���	��8�4����(�NA�\���y13�S"\�Rk�b�����Xu�:�e��k���Mײ+BQx�<�4Ģ����z��Ew>��?�����)�F��
Q��k��e\��$��d����F�ǢK�����v߳_�i�c�~o�.f�U�œ�Nf.����_���P
�%��v�<�v����4+&��V�v珙��̳츝��E)��@����r�c�V�*�7�p9�~���^�w��;x��6jH>��{���m�R.H�+����V`w &��2���7�u�o����1}�u/8K�4���۩�z�B���ӂ������6Q�<��u�#�M<(~,`�C1 �����T�c(�C|��2Tx�*�$~�:���؈|�R�~����^�{P�y �W�W���8OK���Z��v~9����^=�k�qmJ��,�_�
x�+@��X�zpSN�h�����N���v%�~�S_Z����l[07����	�ҹ�3��0�@�Х�zG���ZG^�s8H��s %�����G�Cr&�V�&-��9uvQ���.�w���e� ���5��-.٠u�+�)yx
��NC���c��FD�Ip����@4�����[�:\�-��� j������,S�c���"��Q��THK��{�2�[,ݾ6$��e�Oy�*�8>��5�a���V��S0��8q<��L<���"�3���Ȏ�=�����a;��ɷl0�@�!��1W=�nB�|�����y$�o�e�[�*��9
�ۓ���v�����D\��1A�(T���_C8��ǣnk�Q�����z�6 �n��%����c���E �f��o��[)�;�<ƠX�%�j�}�x��
�mWc��w����-��S[��Ϙp�H�.Xe��3�@�.��F�����HCc���*�n�Z�t�%.��᭣�Zya��ae��q�5]�$l�F��&��⨛�I,�E-��\�cbX����o���S���?�QN���Ժ�ks�FHRl�j���Y��a���+��<�z`�-�3j�ghy_��Q>+�PgQ��vI_��b�G�u>:�����W�9S'}��L;���u~��,t&:�Czh��A��?����龜����옸��EM��>P�U����	���%��6x�uN�c;@=�
F[��1��l����2��m,�����Zz��ޞ_n��J������߂���	j���NC�b:%3>��nH'<�z��_a�����n�J�������3��z�����NJ������v���a�V��!��(����N.�ܧR_@����ur�]K�Հ�N,��N/�i����C#�ZgL($)9RWH�le���z������'�����J�B���z�ݍ1p�N�c�����Y}ݣ���K+�xj-Q���� �)`3d^���LD���^{Ę�
Ÿ6�!~m������Pl����D��聕8$���<ӳ뒝�P�����C� -wo�p��� 1P��waq@PS��ߺǪ�-Z�e�{���:��=��ۀև���+\�1 R;i ���"6������"�/�!�WAB��؂û�����pk��<+��x����h�mI�+a_�6KG���͓����]m�bd��҃wL�4�
P�v�ߎ�M\?I۬�ߥ�����)��K�k&^c�om��$8���x��L���5$.P٬	�0����H���	_��/f3ҼU�+���	��	��ՖM��񣅹x.������Ā˩<Q�7�6�k�,��-m*������C�!Է�~�0��AsKDJ����!���֝�)��_�P?��_�����g7FH����}m�2�)�I,w���v��݇+^�˱C��9Zq^1zQ,-����)B�>��U����"D3�x��C����_�������m�S��K�������h�aQ���ߝ.�����s`wu��aٔI^V��r@��P�{hDw��ni��7C%��Vϵ7���f\z��� #}���&�*h�k%�o���kR�\��i�
c�i��)��Wzw>��2�AuXg����i)�B3�(���~��a���Dǳs�]��"�跎U<p$g��˃!��Ѿܳ�G�.�=Ui��@|�̜>i�tB�s���5J��l
_}���rE�&�Zh��'��	'o�E�I#C�;��;$��|wY��V�?��c�8=���My-ˋ��Ňb��r(�������
�2��2�����r����wg"�d��D�Z�<x^�W5����i�^�'�~��]�ܯ�a�-4gVn�k䪧)���4��[�4���
�m}:��O+��6N I�꒸zǑ����A:� ӕ���A�]��#{5��AU��������mA0q�ˑ"�Db[7f������L���gMĨ6� ��	>�&����	d�'j�G�P�Y�uŞ9�X0���LjP��O�`F�#-��9���ZOB��]��qχQW�a�h�>%�w�x����0�?]��B��NB׳2�jeo|fWج��$m�zL8�8���傹�]��'�ý��|���{��~	�3��9q�sH^��1D)�	�b_V/�5��{�L/�B��O���u�����	�a��D|�ޱǉ�[UW����.=3������YY�֨��D
r7��߁�__a%cup�(�?Q���v����%�5�v�[5�VR�%���w���]�����������g�Z��r������B����Qz'�g�gәF����&k������[��+������+�NV8�%�+8;R��h�>�ޢ=m�KK����Jĸ��Z�.BJ%��U�vj/��^�Ul���s8G����ܦ3�c��@�^/:-\��k5�{.��C��rʩ�֬�/���ؓ�������(��{�����L#�WLe��o��#��3�Qc��Ӕ�$|3����Ck�ˏ�z��woGu/�{�͉@XB���חS��d�lr{u2�0.݀� ����#�=e���6�u��t�?��^r��ׅ.hOJ*��v�Q�a��!������\���Z���zr�=C�ϋ�8��J���L��$mK�	�M��u�Kq�
���r��?�/١+��V5��BOW!����u�!��=�j	"lҁ���`�/����)���Wf+�j}4��(,)怤zQ�;�a��� 6a��7R�"7�����z]`��gϦڥ2��#�K2��R8�,Hb�b~ 8�,��2k�+�ئ�ү����x}˒�����j���oy�h�j��\z�i���*�����+��I�<Qh�l�n,�q"�)�h�y�b+�~-v)X�v��(+&���U�މ$,z��˖�rM3gֲw�I/�
��NN����n��-%h]jah��L�.�rl�5�@\[��B�0���޳�?YvӘ3@��ϛ�1�=^c�w��O�~��Z6��H��	�]5�T ^�J�b9��o�0p��/{�!��R���Æ�:��9�����r%�h�_�2!C����.��aNw�o�8|P�,Q�-�W�����`�e��OU<��<zE �.����1�D��N������� N �:K�d-J���s�X�ǩY�R���<7�>>`~jݬ �;<C����߳��������@V�Cw�D�� �i�ɉuA���>�_pY����n0ѱ��dK���zg��|�G�gg�%������瀢:����C�h46��wPa�sML���.C��oQy�ޤ�lmBF�X��o�+��D���y���G�2Y |�k����w����"/8���`#z�1��E:?�.��]v-���ߔ���s��v���w4�<�eWg�?�OG����M�*D��	�	�X��n<uL�E7�eJ�0���L��̣E��]!7bQ{��D�@��k��)����u� ^!�J ��{`e�&�צjPHƄ`�� ���ek�Tr"c�Z:Y9p�������ο�D�|	BC���[mת�%�Q<l�.1�	���	��=jZ����� !����������p%V��Ȃ{2L�W� ����w @�e�0�Ճ'�  !����Hl� }%��V-Μ�K�dM��r�jxj]�Y��!�� ��a�y��}���<���{G�8�gN�����㗘��mA�oN���W�R>^V���c��Nʊ�v�Ʃ�W�� [��p�o[�9Xԝ�4d�$ߗ2;���K?�#U"?��É�h�& �!�3yh�t��'Jb�3�����r�3�]��� ƽW	?W���F�/���Dw���y�f����7�R��W�X�����V�i˦p��4�)5Z_\��O;`�n?��M8�2�#C��j�|'2�$�L�$A��/�\���hMkܛKe����9�>w���t:���PQ���Ć�9t�5�c��8��x4D��]���>Ϛ�SnepK�n� c�T2q�&RA�au����;㟚�wm�#냸��5�Q'D��/L����h�����G��c���j��<H^�����ۛ�D�,ub���v#PE�\�IN�� �C�?ﲨ�M��2���������Mg�z�j�'Qv�X�C�$��b2f�r�voX�P�q�x #:Y>����7*Ȝ�k��9�Z(g�k�,*��n�I�ټ�cT%+�8��$SߖbX{*�'n޽�p�, O��������W�h��I
5��cH�	�leo�Ff�>�����'� �M���e~P��G�2��1�I6���N���]6.5�s�Er���W�I�t�B�+�?�}�N�'�	R�<���go���;A���q&N��t�p�	.ţKHjhV6����S5��6Q6{=4� p.O��U�H�����J�>ݡ+���/�p�W��8_�žl������`�'�f���ζ�)�u]��A@]��Y� .+@�����q�Չˊ8F�V(��$��
P��=?�&��N�|��
=����ey��*��3��|��mrl�<ɝ�����9���N��J?����X�H�m�L�̬��l�/�)ܖ�nTÑ��+���ly��ﶤ��o4����oe}s��]O�9�ԧ��M��L���A�{jм87`v�U;qY�V�S��B��wN�
p�2��]-oD5}eUߺ�[��~W~H+�:A�i.����N�b5˺��Vf� ��X5�+?�U~�x�4Nw��[��Åμ���n^�I��0��-��^Sצ��?5�R���9@HH���2ܠ/:����K�=u߲�����ŰgZm�d؞��@Q\�@���
�v�I��[(F���@L�AC����z�J&�z�#-�f�<�U$���C���u]�������M|<O�@jLH��J�'��>S������U�$��N�?K�L��Y?�-�:x�<�^�` ���sb�H86$�`�=o�D��D,�����=t��S��[�3�x{1I�s^�.����Q��=QI�q���0=Π2O~ȃ�v;[2Yҳ�b׎ȀF�?'x&�EH:�<j<�:�u����0�8�L�G�ηؘ0V�=M��<�c�5^�C~S�G���v�_���+Z�����h�p�Ŗxg4\�r��~4%G؛�g��{���ng����m�I����i	h=�T��m�=ώCR�5�3q��!On��v衤l���]����W"�WC�E ̾��Z�=:������g��V�m��x��]��!���M��"�z$�!�qג�3u-����}�kC�va�=V�泽�Ь�,�����S/>�9zj��\��nGTd��4�?^������	�;�=�nri�ə��I㧐�S�Bu��(��[�?[WW0"��2A����I`��sһ'��H� ��svt=*[�W�V�)��(�[i���@E������~U�H�Ʀ���4���Q	Zƃ_�2(uّ�}����Zٶ�ƇP,�*���}-�-H��g�6��oL��DG;�W y3z]}X�Q�Au@��+[�E��Պ�'����.|`\F�ߧ<���gHI,]`�_5�&5T*	y.�`�@�pk�QC`�'���g��%`��	���y��*��Q5�Ŭ�O��"��\5�}�O�LZ���/��R�<Ǚ�����Y���&�����3S���QK�R.e#�u�ǽ��Dq���T,x�s���q11����f�]�K��Z4���}$��ɋdPd�	�}�`}�b-K�tW�o�w����H ��ߌw�֨`�(�9k�R�^N�����F�KRj�T�>�L���rn��F�g�q���ގD�O=j�TZ~3�3�="/����N�x5��������jj�@��("�T�"�;bA�Ҥ�*���(���B�J tE��4�I �5@���;��{o�;��u֚kι��guA���:
���[9ILay����Y�e��~�x���� �݀�B��lxE��
;\�tV0��|d����JF;,N#���#�k���?I<�\�72�5�+,�UX����lW�LKvҩ���*�eC��g���Tf ��Z���|����5�z����l8\Y$o��D��C7:��P����V�b�d.}�,�	/�啿�t8�����3` kTR��|>8�տ5��ok���~^@*-����{��P�n�km�}��*TM���>m��>��r�B����V��E]�\Q�����E@DX�
@ح�����U��^�sBo���� ��Ҥ�b��[F�L���0Li�9}�T�#�,Y�0��T*1�ߪ���S*����7G��Qe��*<�*�b8�� �7�4n+��dOU��	�QȾ�K��#�����초�J¢��t�����#3�K�b�j"R*/d�����<�_y{��%\K�`.&�*� �4c/VUA��B��U%����;�f�=g��1��fթ�ˠRl�␆�V�VG���v�� Iqm�r���y���W!"c�3��6����}V5����H�E��&�bbc��~�{���Mfz��3S2��qo�Y��rNf3Kvro�	�����em�!,;����f&н�>A���aM����(���}%ܨK^�hL8��'r�������i��
�m*��#�ި�xs
J>�b��џC�@�(`���*0C$���M�c�N��d�72櫵�o�/�ha�d$�������R��VX�*˜a�S�m1���i�%r�aV:����]y�f��op%��P����"�<P�͸�?P�>����kl��[7�&f�O����4c�����O�,r��wk�%.��$�eB�ŀ�'����O���7�{,��t7��fÝ�����Oob�|%p7��%���=[5�~��1&�i������A�?�X��!_+�'���Co��6̖ȷ6���o�B���^�6
��>�_��48L�`]u6j�4����>91M�D�I��M<�It�w]0k�j9rf�D��v*¥�DSlM��T9�E�}�I��(OY	�n�J�N5����q�7�'N%����0�Z���:�9r���+b�3x�D.��<����G��:7=t{���.ѹ��	��,���h��YҺ��,��&l���J�����r0��̮�N���"�>���Y6�x���i�ƙPAl���g�jA~�ĄK(�z5��'S,~a�ɢ��/[?Sizf"���ֺ\�<U�:�I<�cP��6:"����+�x^7�[�TafM���V��)����g��R6��#v2;�m1f�E����9������2�r�Na���?N_?�q�����݀V`�o�E�W�943�(���s�ns�Z��z>FB#/�efg�7���A(���Pb�X��.���K�÷�N�??H�"�����9�k����+Z�������ŘE:ঌ�y���G�$ۤ�ڋ]<Y�c���T�4��vP#��!�Ib{��Q۱�	�7��u7x�-u_i���q��9�4N���$`�E�ǟ��wZ�M�L�� ��1� #Py���b�М��Li�z���у�-j������[���5d[탵���ӥ5 ���w 3:�%?s��O��C�x�j�E����'~"�^Ti��H��7]<5����Җm'}m�=��N�,HU�2��*`o�Ԧ��:��Ur��hgw}��͍�!'F4qrnI2`��,���{CS,+W1!b�8��(*�	 �r�����6�x,c)sz�Q����>�,8X����f����Rk <�]po�����u;V�X?��S;���߯��� -t�g�?D�#pyIm*�14�W=�%����:��B�
�fꧢ�B�WO~��d�_1��:�CDe�$X�F(*�c	�)ڃ�,A�]�����RR^�6��䈟BO.�t�=)���'��H�Dj�eK}Ǧ!}\�YX�qq�K��̢:��30����x�
�䇻)/��$[o%��YV�w96�g����ES�os&~a���2�.9&�f���u��I����o���/�E���o��;�n0��D]�v��"G�'�ceKp����g� �\��Ԭ��}O�$����R�ud�Bo��m'��@Z��p>m�tI��:�/k\@����~����,�`��i��l�%�q&ދ�87黊>�)�5��G�!i�S��1h%��Ƴ�/�� ��dY��v�|�d7;\Us��l�����f%F>Ӕ1{	1���9�C]��mh��BqӲ�����7ַ�������(��@B��U�|���{�ؠ"뫺�TBj������WS#���3��Df���E'���O�f�N
1t�K�RG���G�t��6�O�V�L�o" q��q���0�Woѭ�{�D��k
W��Ơ��?RY��*�
;����>M�e��s�-�lc���s�1V��3~�̫��o�����r�"���N�i��q�����NoB�P+�Qof.�
`"Zش�?�w]X�eE���`D`��r)`������j��)V�/+���>t�>Qi��L���P���J4������)������12�[Z{n�	�B����;�K��"�<kۺ���\o	�f���� ��4=���q����o�=��<����j�S��	��}���̡M;��q�����]ٖX��Jgk��05I`ZykH�[�=��������ɭW��g�vb�	=K=�aq#����zY��G+�sù�1C���O#��t^b��j�	�����rBw��5��/�}:�X�Wl��E����J��\��Y��F4��Z�'V\%���y�J�L��W$�-���y����ܝL/2/g�5[�;���¥f;g�43�'�Y�̵�����ɎN�#�jR-|�-)o]��!�E�'��D��D�0���1��UҫR�XD�}e��68�����Hm�O �}��o�~{�L��l��✢�����-��i�T���cei)���[���?�1�{�4v���ӫ��Z�|� 8���絻�mC��|}f����g/D7{��H��۟O^^��E|Oemym��D�A&�A�oy}-N]�?͛OZ��jZ�n޺EF�!�|�9�X_�~Z]���MzEq�}~ƭr�Lb���㇯����=��H��UI�a�8�S��p�E��e5�g,YǮ�Ȧu� ���~�?��{'d�f]�ik�%����Y	��W���ZՉ(�{��0OCYD��8 �y��Y��9n]��L�
3��+�6�)���	a�m����>y>^`��qKͳ�q���`��䐩���<��Dh���;��n�e�ن�òY}7Eo��e�Y��VG�|=b<��:��g �0t�"��E��E��F�X�8�f�~�d/FN��4au��.ax���}�+W1�vO�@ȵ����q�h�4��;�o��锪H�0�2%ɒ��$4�	�y�fG\:7�U�����r6����t�i���w�*~�H	�V�/r ��w�p������P�d�ݾ���p������r�O��dפ��uӖߊ�O�������5e��fB�p��	���"�m"�F�y��*�/m<��fI*0"�Ts�寑��B�`�1�P�KXy�}���P�0�O#E0�/�ˡ.��g� �q�P�'�9�+����/��侱q��5�.���%
�1�� cQ�^�����+m�����!!Bh���Vl��6ǁ�,w�����Ŭ�,�m�nc�-0i�3|bZ.��n�&^S�'=������2*�bF�ҙ�S��X'�Y��[�,��h�f�cf����Yz�%��ys[�W��B2�6�0*��-�_<�8e�̢!D�M� Mq�H�i&�d�Z���]�pF�O�E�
�:��EN�����%ͩ^�Q� ���N��;};�U�D@�2���9�;�8%ɼ>i�.����*v��X+l�r�-7^n���1�V��֯d%J�59��WN�j$N	��+%R��oz�%6b�_�O����o(��L��^oKB��[������&@�o��T�֒P��%���B0���d|w
��
�Sl��$�������};t�f�jS֨b?�A�c�ڲJvV�D?�F	Ȕ�<H��m��&=�]~�v�ݽ ?�Ǵ������Ȇu��<ƺLB;��>�Q��I�S࿸rҩ��e2�=��B�0![#�͘/���WY1���r�C�[iD�$��Q?�B�ڹ�j�P>d�Џm���B�O+y�w%�.���K��馮��$s�G	�l�{��� g׾�V�^�i��d/5g��|T�w~�b��W7S�� ��	7���c�}�2����/�X�G系t��1;x'7�
r=�N���U}�����G��l��#��uC#7r��㱳�U�6:��s��|�2��ou넺 |��[��-W-�)�&�\�N	~ba�/"V(T�jQ)r_�*�s�T�QXE�J�v�DdJ�E9oy&��)�� �����l��H!1#M�P��tr>Њ�295�T2���ϯ��r\�����(���u�o���ټRhrT�Ќ������ �YF���"5L�ɵi�1�uH2tB���aL4��5����tk
'�q��w n�%���?��}�t��˶y��8I�H���_��ۼcip���~d�li�M�����'' �CD#)%{��
��>*?O�	H0��v;�Te1L"È�.ek�P�y��_j�Pv�`]ϒ���WM1�?\	�ufgb �`J臇d��q���vqP�K�P�hOF综�!}�K�(�m,�M��k�Mgڨ|��m�(i���Ϸ����R_����j����	޾�,�^J}�������5���U�:�+�M�k��A�5��~����@j6rß�L$�16�o��E˾���k�	Q]���E3l��닐�N�Sm�O���U?Y=1�-��Kt�V��c�4KX}�护��J1��sPg7�j����n�g�1?��N<����ֶiM��}0&1�q�6(~Jd����ط����9��)��8Ó�g8n\�N�#3�nqa��[K�V��vXhA��%��FK'u�ej_�
گ"k��+@�-ق]0��;�.��*NLB���SR�T#�WÃ<8�n���/��_�5]t���;�4
9�r���<�fV�#�����aH���ǔv��i�}ָ��0nM��U^�rVf�"DT��ĂqpV�_z��^��%���ʕ���ɽ;��	'��1ϗ�6@��F����ń>���GnѤ�p�!:\�d7��rT�/���ҤϨֵ�z��ࢄ#�دԓa�j�[�yfgW�xV�|N7��� ���h�a�a�$4)i<����}gj>��Z�&�՜Se?A�h!}X}�=�0��Y��(,.V%ǒ��R�[^�՛7p��%��r�������,���w�e?�ce�e��&�p��j�̰g�y�#vW�u"3�X�/r�pc�z}������Svsd c����U�ԫ����9_%Ϛ��|��RkQ�����( �72��Ez�|�_U���������F�M�}8��Ԍ��8�'���}mb�?4k���	hf��3ϣ���b�
uI���x�G���=��.�d����uAw�ȑ	n2��������O�r��0�oago��Z�u�*޼�K=�G�@���k�a1'}�'�<��E�w�z"`m�ˀp�V��Dq�ʝK��3��b*Y��)����,~*�o �O���In�f9�e��#䈓zݚ�~fw2E��x<��������g��_ݯ�F���U/+�RQ~S��hB�F2�W�K�#r�������S <�Ub�$d���l�Ve;��a��+���M��l�;�｡O�8�����������������ϧ;7�He��=gdv������C[�DDv1k_P��
d`�W0�����$8<,H���i��[{��b�M�k��j��4c�u��2�ך�̐7��?^Hª��<�w�,���Cf׏����(�m�\Č튂L~����\L�W��X�@G��hx�[|3(Y_����z�ȌNd�*��ܐ��.S�4R�8�q�}��ܸ���3�,w�T��?����� %g�%6����X/�v����%&7����K�g|��EN9D�H��i���9
�N����~+��
�0��J�Ӟ+�+���.i���NG§SQu#ē���2ua[Ȳ��yʐa%\���xiI`�1~P4:���̓J�F��Ϛׅ�٫M�m�n:��/N>�>ўJ�?a�t�؆�Ψ(@}�	�a�i���}d��;�U��O<�V���9W��䶊��LJ�i�1je��˓G��QE�ޱ"c|w��W����b���>"]h=��q�\��j����?�5k�Y�=>�ɶܳ8�����S��e����w�2����X�S*2��_��+4E_���w �p�\�t*��GP�V`<�и�$D
�p�i/�&��a$��BP�K���W۳U��ޓ䈚Q[��9�߮�L���f���rB�ēq��<��8[�MG����@�!r�W���pV}dn����D�yS���s�T,�d���N�§ᨀ>�O���ra�|����11�e��=��k��*˱�{2�`qC�vgP�� ��sw���X�ɾe�B
�nX���b��nv�¬}����[1K����>g�[Q�쇯y�z%�#��.�?bb���P��C��E~���br��cE��di��*ٛ�Ќ�i Z=7WY��]Ɲ��j�0��5 M�Jq�t.)%�H�;O��y9>Vh	5[v�U3J�b!\Mމ8k/6��ء[1��%�B��ֶ|x��8�\_�T���mx�����|Cv�D�c.\Y�H�^īkW�2��T�sI�tr�O&Ja2ή���7���鏉��y��$/׌��{�s�}\�W��-p�	��v?W�W���Ͱ_�j0�+5{X;��X�UG��� ��-p"%B%]����-̋w|�2�`��<j�pF�+�֕s_����Ņ ���ľ�D?�؀X����y�2�*w4y��`S���!�fߨ��bb��	�Թ��݁j&��yj�2TZ�s>�E%̨��Փn-ċa����*�B�=��=��P\�1�orP�è�m!�9A�	ΰY .���㯉�X�*:�̛�����Q�DE����/�[��-�WȓW�$��c)@ �a�T�Rp+�CLˎa�O0o^\T)#����CF��X���+E5G�����SS�I&*���Cw��;W #�i¥��6!\0ܹZ�N���$���Ơ��*�|�3���5�R�r��t�@(���}��ɠ?������}Bش��FE *N��m�5ZF���Ci�6�*���� �M�P�O6�-W%W2�"fb�\u�| ��;w�u��g�2�]��Y�
P�T�Ҙ�֒����n��jb넴[~�ޞ�x<J7�T{�RHq7
C�y<D<���"������ç�N�����أl�D��QLB����%ꂪ���n�0�6�j��_l*ԇ0�*��e��I=����M,V�:����U�\8Q��kL��_�����F^��{����7�L�p��b�q�$o_E�"���y�Z��E��x�yb#7_��mn�W�]�����9���b��~���,п=�L]2ޱ�����%��',���J�V�F�r�%1L5|C��g�,�v��o��G��bCjfJ�x��}n�tkH�Z�p��u<e"�#�E_SɭA�ܓ։�N)���,pz�;�h���]�(�?������0�����B�te�
1���s�豓��"�*�z@֖|UTҵL�0_��)���əqI#��_P�S��N[��ҩ�fG���|9�^M�����P2g��V�e�tw�dn�I�2��M��9��/Sw��G<�>�X�"|��7���wVleW��cx�*f���r¶yf��$��=���;5��:�4����A������_��%2/Y�I!/k���g/4���?i9�8���jSA��<��NxAU�����\v���o|)�j���`/^��e�k���_�;|;ґ�h�0ߪ
���z��^�y~��� �J0xqQ�W�380���B��@��<R�2�8N���2R
5 0��uab��zz�5S�8Z�I5P����CnUǈ`��b�]<��@~�Z�ŷ[z��p�N���˾�$�O�E�/��|�?���I��ɹ�P�7�A^Mp��y��9��d�P6��4�9���.��įx���ǻ]C�Q�q[{��!���IR��)�P��K�x~�%�oę[,c�����T3hWa}�;����#�Igڹl|���H�ߏ�ɵ�
y���Ќх{�ฌ��F��kB+3l���>�#J��~��<�j�8BhA6<mKHˣr����S��	��Ҭ[�s�p�HB��iN�@�3~ь^h���k�+�l�[ڡ?y�q��EK%��_a�a@	�`C)�}4�P�W@sP6�@���.����0!�4�ui�@�r��m�j?���>oaaЭ���
P�K��H�]�*����$Nb<��ל;���S)fM;�l�YDCʢEޚ�F�y��T3{O�|5
���]�x�Y���e�奇t��;#q0yO4W� �t�ldkO@����+g�����ch���xa���� ���7;J�sl�x���_�m�
�Ҭ�d�:��)7�a\bO��F�2�w�:yX��H���r�������$�U�u��Do���d���ñؽ�z�F��64���6^G%U��6I��0�~���t$~��#m�݌�*�3�0ް�B!G���~��z���%.`5n9S����lQ[Z�F.�{��^�{#G�/t�c��҃o@���|-�ݚ��l" ��O�5L� ���0�QS�HQ�I�p��Ϫ�خ�Fp!�D!ZNŰ����{cR�=�]cvv�w�n{��);>��<V�3f��
h��w�}��s;�;��6&�2�\�J^Q�Avr�\m�y��{�N��g[?l��ʎ�x�:�7�_���ۥ�Ќq�k��K�Ϯ�?|���ɷ`��#l��ù��"��n[�T��'�`xy�r���,������W���ssv?:g��E�A+���I��������Z������r�Xw��f�1.I�؄Hμ�u����p4Ai!Yi!�1��]���Z��������u�������9� ���1s�ʿ��-rv��S���*껅����%�3ܺf����d������w�n��ùӥ�6v����иפ��v(+WJ���8�-x��B�6�RG�X���Ќ=4&Ո�pv�]�򗻊����R0���.U��01s�XG�������py��/A �t�.�k0=���5MI:H��0�~i�Њ���y��x/n6�ܰ\���W/˝aͿ��x�g��Wz���% ����z�)�@�ӿmg5�j$�٦� W����G�Pʚ<�P���.˲:nq7AX5c�,��ks�	32J��m�Dp|���[reEo|~�h����Ѹ��C��0��{@r�3�us�ސ"�6���G��R�k��C�ΰ�'>�j῏���6��Mx�v����ȟ!�1��@K����RHЦN��]�/7ļЅ�k�2�bgWU^���ԡ�o�+��t|�0�!���[@U��d��I�X�[�s���A�7ee��݈�9�gOU<��;����Ƃ����c��[��2��x-���K�J�zt���e���m dF�8v�O�TR6�đ:��;�1�ϔU/7�B�o�9X0�E������n��lL��B�(-{2�c���%��@�W��10Ψ���^kvy�q�E�.|���ؤoRh�Y�e)ww1Ŕ�˜�S�J�f�kRY�@^��)�MSZ����H�+���$����:*���d1�R�Do��q,��kE�����@I�o��D:����!: w4У�� �E3G�ۮ�1�.e��Kh��`���a��S��\�4�8T��;��<����<����>��T��ާI3X��Q{Q�xT�#}#��\�!��w�C��/y���Y�E�u�U~ä����n�6��ֹW{==�c��pBQ0���1xo�+g����P��L�����}�+�^�.��taey}�;����-�7^�{ߌ$�Vi`0�z�ˇ���[H�m�7�>�I�D�I��ҷ��%r�6-�w+����!f
��2���1<+������e�Y��� �][����K�Wjb�� �Z�Z6x�9����/����2��K��6mM����Fș{<E��̂���K����vЩª��B�.T���TU�m�o����@�s��t9{l�EJH}�݇���n�&f#PP^��F�����ݓ���m~ ױ�@X-?�8u�<j:h�7ӡ���=#1!ִ������r���ϰ �[�ʩ���L��e��KP�E��:����uvЫtb��q���:��'�hYL�!-�X�({Z� /��y8S)�����8jVwB١v/��j5����b�(��tD~	��e\�z����B����jYF����j9����<����#�!%d�İ���+�r�:V���ހlf3
F̥�j����� #��@{�9����lj�fŒRf9�Z����q�!��!��6!]�wb@�vA��4��Q�@�G�!��z�@�g�P(��gK�v"�<V�������˅�̍���R7_��X�;>��L�D�
*�S������.	p9o�+V5��{�&Y�@�|�.��V�`-��#����B��0x��AH0w[I���?��%/,t߫��>�o��Jf���,�Y��	��!�gH�d1{@%j ~�'� ��N=J��,��]}���Q�hzupo��mGJ�֚6.���e!J�&5YS�����4�,c�tSK�Z��^m��%Ԍ:�-c&���|���N	�S�O�~���Wv�^�(R���y�3���l`���y.wNy��ϥ��*��s�G��I+��>2��ܝ���},�?���_oX_P�Sq��(/���	���J;�i22�h.���FMR�]&���*U�T�T�J�퀴-W��W�����e|m�̤7t���mE6(�SRd+lb�3NRk�\E�j/V`4}���yulp�|���WA�mK�;k)�����"&� �l��,�f�t����� ^�s�PDp�D	��T`hM�&mp���n�F��#����!s�j%%�����Eڪ1��%���ֆT#����Ȇ>�X.�S,6�lI�q<�o�2Xz�(���
�g�`���<�
��/5�[y�B�8o9c�w�˝�\�\"�;�Kr�-�ՙ+5d�ac���{�U`���jþ)g��x���J�&�<Pe��8�Uցݿ�?�G���,�/��^��J�O��n:�/r�]jd!��_���9��
�H���W[�!+��E�/�g:΄������C��m?���ؗ�ˌ�l�W�6�j�q5|�����Zu���P�هe&�j���dk�K�O9f�W�������!KX�J��4��{9&w~�,��*����H�[Xz�����)��@ޗ��-��65E���L�ӛi8c�iA�~@�����;jl��|f%_t	�+8�����w��s�WF ��kw0�.�Y�߻1!�m6��7fS�Ў"�>����:E�[\���|��-ēf�f6R�R}���ͷ�F�QE��A|�Y"w��O-pN>�gHm�;��40��x�Ӆ�G6'���	٭�c���6G�fv#ͮ,�_�Ϻ�M���0����/� h�ΙJU7�,���Ak�������<�Ut!u�P5�v|M���w�hϽ�ߓ�E�܀ ���{�>����'�]��G;鬲�]_)*�E\;�5��9|@�=sѰ�m<�ou���;�j��#���Z�>�]��2��`:z�ײ�W�����:�d��T�n 8�EE^F��^�j��� ' �p���|�3����>z���?�g�{vr��g�����}$Zη�N��~��oy�}�-{��QC�_�;Ě�Bhso	�Kz򊘦������]2`Z�g��Ϊ�:����ɐ断,��;���yoDZN�h��>�X��ԐHYz)�zBҸ�0��m1�.Tŵ�O}D�dK�������^4��NC��X�1��[4��ˀ�y��m�憌޺xG�?���*�l�?PCC& �i�Q�c��栙Z����*��V�x��%T^�hs���b��پ������,�׀*ѵ���|5 z�� Mz���d�u�Q�,�r��b�ю�
�����i2ސ~n��d�F��_��Fq�=4�U%�xAUf&�#�'��TV�[y[��ˋ_`宜!]�F�?گ�W��j��Id�&Ot��}��ꂈjM�<ŖGC[@����K �A@?v��r�bYh��Ddo�m�ktOet�m+W'j��$y��uSh[~���_���9����𰢱���U�^D�8�T�MbdJuY͍��eK@\\p�anN��x"�y�HJ�Q���5�SS���Z�?�ɗ��^y�<����29���!��Aࢋ�M��C�J�3��)"��>�8���*j��oI.�q�uβMs�3�F ��3��[OZ�5	5b�Wɾ12�
CC{ �a�bK�{a"yo3���/����?[��o�[���c<E�~��)�QΡ}��w��>2��@���0�+����s��e"
)������8N��FC�,,��]:~�l(Y|�����/|5Nf��Z��Î<��gR����z[e�k��0I�Ղ��X�بʇ�, +�q2��������R��kB9������Ϊ\b���Dʺh���E�A�Ke�{'אw�Y�Wߝ������׋��cs�����22uaZ���ں�З~	���v�5|�T#~�M�+���F�M��^����[[����A�f�����֝Ҙ�¹�G��֝���
���0ghxJbڏ"�n�u
�� g�eV��&>}a☛�k=(B��z���#}�r��p]�9����nm��d��A��q��V�<=B0���	mA�����b���T���XhŦ����P�Q��g���d;�e�+tm]M㠑'V�I��V�g�.R@$�˯	�$���V��,�/�d/,���p���ھͷ^-����=$��Ok���XH�H��O֓X0'Sm�֟|��O�Ξ�81�
�.�Ӟ>i(F-�V,Nn����?�c�"�byN(6���2�s`�v��:`�K���Fuӟe�m�A묚E�a��X@GJ�����B��e�E7,��t�T�Ƙ��>�?��d��W�l腫�����=�z�����yEt!�o�GJ���l 	2&~M��c� c0ѩsk9�E��J��M�o���U'ځ��П��J5	�c]C4������
�^�ϩ�����~���v�/�d�4qn�E��O�X�+~E�z	0�3ߋ1l<�7�LI"�:��S+ڟ�!��4��jӽR=Y|�Ӳ,��/�^�o���H�-k�~�y��a�����zZ6�?;��9��ůt��Yfy=���V]�;����>�`�<�U��;�{3�!��w�B�<wu؛�8W��~�����?dεSa(�p2N�4�x�d��������"�� ��Q[��T�}����gH�� �pu�c�aQ\��	τg_=����5�����	̍���h@"�3�F�3�Ը�L+yDrڇ����P��n��9}���EΫ$�(u�����j�{� ��E�}��?s�C_� b��@��7���J����O��R��1#sH>3��=��0�(���>�fq,��13�T �N������� #�'�CJ��&���.���0z��F~��}7ͼ��HE�ײ�Q��i�X`ܙF=�M�vw���B:?���W�P�ذOä�lx��<{�]x%I��H?����z�q�#I��q��U�ш{i�m����#�fC�Uh�W-��~YZ1��ף� �r�I�uDm�����5ts���MfH��ä��/�D�]�N��G��,��>t>&�GiF��D�i��2���p�5��t0ێ)���τn�;�&���#a���0��=a��Y�F�6���(���	��.Ҷ\�\���1��������dc���7諢ǣ����1"��8�̇��v0������!�T
L����-�Qj��o�4�r�F>1��(>���d��`�;��A���2�h9 �8/�s���ڐ�@�-�� ݚ��nj��m���_Q�[R �F'zʹd�U��L�hl4�]��3@(�xܬ���w[~6�/�f@�62B���-:Hi=�XhY���A���WH��>'%�`�Ow���H��ڹ;���yj��ޤ�6��V4ز�Bgo�r�GՉ��
ÀѴB���M��Y(y/{V�:��B������@�J7�-��� [~��G�������Q�i�>a�(�޿��sٙ�����
���A�qb��	�$%�]9�5��R�R�T8�,��	Zđ�����˙R��x�ӯ/��|樳�.we(�,~�<\�ٛ��/~d��$�uF,�I������2��w}gA���f[���Y5��;�|��A{���@�y��"?�^����S�*�	�� �'���L~�[��H�@M�WX���~��Y<7��N]'�Ҷd�	�w���jD�ޘ�)���j_��J�i�ٚ[Gkn4�z"��[X�@~@&�j��i�^~���줕�'��\FBc	�nƈGۂ�1C��N�[1�U�����^h�yf��1��R��e��$�r�+�����LQ�&ѹ��2}�/����*�f[�i"d�M��n�ŭ�d�*t�=��	ԋ�R�/�#��� z+�ӎ�D��ֱ��7	��m�0������� $'�d�=M4�b2��EB��۫����c�	�*�)�E��JE(pA,/�	a����WBb�6Y9��m_��K����U^6GK��u�����ӌ̡�t�#o��˙���SXu�l�WTM�ȭ������ݥ�.>ٹv�n[b?��t��n�xr�K��3������ʽ��K�t��3��ќ5y�Q~��J<�R�����&�#> �^*g�)�R_|v:�W��&1&���K��D�s$9e�}��Gd6�/��R%�cË.,��:!��	����z�������Z���66�b/�8����:�/��SqŻj4��5�`��
��J�@�D��(�(��x�	���m�\�fk��_��a��	��w<����G뼈IG�B��=>?`��̕/�	~~[������Ҕ��/�I�P�q�� �"��$�a�EW$l�s~gh���K��<���e�ئ^Y����[x/���eM;����V�΀8�寧�<w�G�Y$����1{nDL��n���r���b�r��<��kJ�����������6�2�)����*�yT$J^�/��?H8���lH����"��G�����Aѕi��w�����p��ٛ����/ZX�f&J�k�s�yH ���vdc�*�%_�t&�|u���v�Е��eK�tO���J��B�M�hHL:���6�ѡW$��CIF�:q(��]ٹpF�X����G��$˨̀��Fɔ���X�^�ڷ�O���w���|�cl_��u\���M�Zi+�0��9�5�����X�����o;e����`ϐW�w�X`!��8�N�֦.����[9�Vg5�/Sr�����U>=��p�+L��~ӗD�D��������q�ڛfYm�L��3��tBg]دF�N2Ç/o��Yt�'�K��6�+�~aۍA-	��#vQ��G#d"����k~��˳�+[#T>aa�^m̈́�Xh�v���������ѻ���h�Y���oGJ�o�>�8\<�����E���z���:}���y��J��b]]�7t�~j�uGd��j�f"�>����O���S�-���c���7!6W�/�M�M��.{.�Q�b��G���g��� �#��l�0�'o�l`�|Z>�Pz���|��s��T�6����#�u�i��t��9�4��m׌��c'� "z�c=�)�[hQ��M-S���Dӝ��go���5-K �Q�"#3(j���Ȇ��`�O��~bz�z!� ���T)�f�ӄ~��[x|���3�q�x��$а^_����N���o�J0^�V[�������}����8W''M5�g0�'�����1쏞)���I��q���<�w	�0P�SzY��2ޕ�([4�׸�^��n)vᓽ�Z�7�}p�ܶ�ïh�o��Ë�A������w�StfI	�Of�2W��G�j�E[cVsPG�����[J��3�{_�����R>s��ɋ:��eD���sg�)U���s�!˰�#ky����Y��<��~wۦ����y-�s4��s赤�_[�_M�~292>�7��0&��9��f�{�"�듳��L��[�p~n�����ǽ�x�[�W��)J�F�g��m��&�@���R����)�������6��^����ɷ$0{���"��- �/bk��lN����b��X�,�q�SZ{����]�Ǯ��WF�)I�u+�-q4�5ץo٧VF��s��Q���04����D���뇱X*�#9l���i�O���ܚ-<��Z��z4�����s�?ʀFb�8���//��3�,�g���
���.>Y�`�^ a�I��:C[�{��^#�h3O��ŧ�ج��O&�[z�<깾�]#=��l����u�/��[��X���!���!�}�>�)��)�8�Tc�b�����b�(�����A.d{$��|���JaDCf��Ë��3&9k}��\��t���f�}y,42"O&0yC��B�[F���&���K��[I�gYL��_����_�֙�W�9�6�^�s#���<����R7%QD��T���t��Pd�I�����f+�)R1D$;ٷ�dϖ쳐}��3f��<�������_�y�s^�9�y�\!B�v(�Ζ�6�vWK��ԁɞ�
�1�O�wMk\ׅ��4O�Z�/,_(�в��,VR��ϧ��^���O��~����B����#�� k���ɳ��XD>�=�?�rsJ{.)=a7�R���8�X���j�l QC����R)�R ��u�iT�����DXYRT���;�_��F�ޅ�;�������7���\j����U�r|�-�f�#�_w�h	<�f%mRa�+c��SJ�/�����I��}�`��/Q �^���b����J�T�" X֕`^�ew���)[s��:ߖ���/�ǃ�<�vrO����:�� �'����3^Z�1
�E�����mmǂV_6����\��j|���yU���PoC���:�)A�� ����V��)!����$>���5�yWfϾ�c�,>�x]�t��@O���3 �� !��\��2��7S�j�d�Y>��S�D_Es���	���=%u�G��Yo�:������M♜�֖s{���%=?��R��E ĉ]���'���s7�x2`����&Dc�����a�"�$A+�m�]��<Z�}�as�6[h6)\�+�NM'�����\�@ᦕ<��^�T����Pgq��H�Y���/�3me�9��ub����;t1RY�4�{7�����bE,��n/~���!���!�9�#�4�h�����V�#��!\ߡ�ǲ\�&0of:6+�Q���J	b6����U��v�i�������+�)UN�i�\1�vR(��O�.`[E�/�$���s���jȲS{u��ԿQ�Β1���n�CA����|z�O��Ȅ�r�Nq<�L������P� �ݺ��(��u�y%, ij(��g��H�}��0N�l;��3���b�2nh:+� ���W���f~y˅�}�kr;�d�
�� C�ꌸ��f��8�L�~��ވ#��5�zՎk|�9 �Y��4��G�	�-I��BÒ�J�ф�3PU��c����'�$f_�=�.zD�B��a'W^�������v��̔�d���3r��uG&��Bֳh�D8AŒv�7��b�B�Xc��Oh(� �q�zz�_�X�� ��O*80�~4�ҮV[���D2�n�#�gD�|q�< G������.�\>03�Ȩԉp�ǲ�s@'q��Q�3h�����G�6�=�Z*��ʚ8��B��&�4T�;�[�8�м��ͧ���ȱ�c3{�UX�O�m�x�R��/@��{�[4���S������;�摪��G)�/�$�5��J�l⏠T�k�&o���c74���V��罹��U��t
���ૻ��5�IT���d+�ѫ	=�jn]�U�e.�r�2�����%����i�O�����ms� l����?�7ڲ�X�'K�>��W�{)�Dv��)u3P���^�A��Dh �c�����?Z��;����}���r�@y��X�&?ي�
WE��7hrİx����%��S���n����i],0�4X�t��re�i嚫��ָD��ʕX{��95�*�H�Ɛ�h�dO{���^��5�ĳ�����;9Q?�W>��*Ί�l��2��IE�8y:�M��Q�jU��������I�y�<���zX\�b;)�]^�;��b:�|V�%h���@�g={z�}�/�C�c,�����g��Qaw�" e��5{��͛�I��S���B����HɛN%UK4�@�����AO/ru9f"2�ψ2�}g�
��h�n�<l��N<�>�K�I_2X2�J�F�T���@�W�:U�$9ܪ�M��4���y�����U2��	��H�}d[�A�蟾�͹2b�%�.�������!���!�=�P���P��2}>(�ZM�\4@�����}��k�Ϩ���&t�o[����SL�h�%��Q��W)	41���ݳD��%	[〉1�I&:+�O�	�{(��X�33<��`�I8�Yx���R���0
!��pQURĐ��f6%s�h��@R<��b�P���_����;<�1��|��o��^��z�w�F+B����~^�f�'�Qi�����(���o��Wt�"��N�
p�e�\��������u]�v����ɋ;�r��t�{�#��r
b���a<�.ݩƹ&��<LDl���3#�Q�����e�I@veʒb*ǁƏOF��Z�t=�ƥL�_GEs4�k��]H��Ǵ���9ݯ�1	)���}P��9�V�|�`�Pm��vS�#����@�N�!�yH��Oם��7��/� +���㶬|�}p��
�5�WF���mg�J��R6hIH�����8֓����yqu]`D쇚xgD�z�64.AE��,8����3P2�;IX�����;[��:�	̦�@��v?&�~>�vKxD�8����=aA��Cm�� �'����]-ڸE�q���"sA�Z���g��V�cv���O���s{��I?H���'��82�2��~o牍Ev��VwmҥA"�)ԣVJk���Q���g��c�ܐ�B������I��=S�C���@��c������q|��J���z��n��zG�'ڻi=�q{� !^�B�j����՝x�u��ߴϔLp?Q���r���d��;7��n����s����:	�1�	(2�'�E�O�?����7�:��uQG�y&Y@���]��F��+�ю��t'~��f6��SR �[� x���;��x�$[ڝ.��͙��!Y�(ǔؼ��;�,)@V`7�O|�]m�ub�'f�)������'ߙ����� ]�����U�X�����
k�M5�wz�xh8��v(�r�=�p3��W����`]�@��:���KxW�zu����q�@�2����Fj��}���GP�
i#ϴF}l�t�:d�{��� ��PR��/@��ˑC�I˄$w>��"�
��&���xu�������<T���6�~�l\j�����v���������7<�.5f�)��c���/�͸O5��	\y�V����4��5_E@h�W�G��=�ȯ��gc�AP׈��"?��Z2}ZΏ#��4e�td�С@�f3@˒���*в٤?L���?U���s[%���l��\)�˨M��g�&7��*)���t���o:J|����A�D���qj���`L���4&���J+/�9A���`�%�e'`e9*�i���։��NH�\�\�W"�iӬ+΁[@��[�iY}}
;����� ~>����W]z�4�p�2�؄��C�:�����=�W��Zn���,J�]��W�������Tt�v6�#$�.a���/��r:���jպ?"l>{/EL
�AK��\АR���%@��k� PC ?��`e�n�PE�.B;���>*i�G��7����P�@�6�j�A}��;\�xq�r�_*MW]v�j�ȟ�g	fF��?��|L����ߠ �.���5���V4�^��u$N�MM(I@>q(�x�d�P<Ю�ϛ�so�U�ۖM���l�qM_e	�g�XL��q�*H,���=��ϣ.���B���:T-���<�pj�*D x^�79�χ�ε��W7�k_Z��n�1$�pRjS$�� ��oau�w��P�|����n���*��ó�8����B�4��i1�{���o�B��}~�Wܥ���������**�6�	�o�a�9,�zZu8�:F�u:���>h����]�\��O�Yih�4RZ���S���S��,ޘ�/���>,|�6@��ɋ�c�p����=�x=�;@�����3�|�=3��랠V��{���������0
n�x�
��
�e�"[_�������%���ߢ*-l,��@u�������(�=�2�a����[��6vhxh�P��p�q��CRC�2��#7DN���E�QV��o�����x����l�C�W���"d���@�9�ㆁA3�2��4���y^��@tG��H��'���C��@#}6�T2jt�mh�МS�O!C��޷�,��ing[`k��Gj~/�	�[�$Xs�|��x)��c=�GB$*�hX��ѱ������lE�����q�@�b�wVs�^O����"P�}A�)��3��;Ra9���w��1ͷ�T=��A����n�j����\e���Es�
�ҽ>��6���?�0�p�?�6�>�j¸�r�H���S��j��rF���@`�77���V�l�-�+h�إWdj���6� ���a�%� �%�i1�$��nJ�',OO ۺv�� 6� ��#�_�{F���ފ��y`��fOA�ٔ���Cf����fx�,�Xu��)���v� ֍��z�x��̙�[��[��VwS�_"�i/$5PG����7�Ҋ�P����f@ӀŦ�C�P�����T�҇����Y��)%��-�˵���v��R.�O�a�ˆg�tj��DJ}H0Nk</NI9�a���'�h�6@�a��xQ���)�$^���
��:�?��[�!0�����\Qg4�CX�
���x���
��y
����p�o�$ӻ��0�ة��p{/3A��������.����--��w��u'Bu*��5Җ�m�� }��kio�]��ʺ~��0U/r��(2\pPzA|������){������<��d/!S�tС�Cm���$
���ܣ���!v��f�#Ûo����M�����e�4�\{ �A�)�����}�P���T! �9��J���OEG�ʭv�;ϳ��k'5�9�1�+�D�a��C���&�	4j$|b\IK�8���y�Ԅ���)t׭��!R�7t�c��O51o�l ����3߻�P����G�42|�ye3��@�1ʽb���(vK5	m~[Oc�"٨���[#��D*J �"�h$��Q��l� �U
��Khxp�'��4��T�{�v�o�X@��Z1�F5��l{���	�g�3a���k��C>��5�Ng���&��i����ģ����+�@�GH�Ym��jt�$��*u'��t�> ��h��m^|JשCٽ n�*#G�\_X���ɝ�(�8O�Q���`�Q�X�a���|�-q:�ku(��������~���/,��=j����Q��Ts�L�aef��d�;Xל�g��yE��+�SE�sV���do`=#u[l{��r�~6?�u��`�8L�>}M;��7��_�Q��y51�?qX���*��A�B����!�S܁�v!�jx�h�m�2�;�l��x ^ �6| 9����x6�p�����@�R�٢�w�:Ō{�pK���4�ԂO����R��ii?o�;�L��CxO���o(��S��H��&AǱg�3�w��eMI�O	�k��$���O�I#���f�	�s3�NU���3a�"
�sr�qU�oKܴZ4s����_��6��n�c!����������4�V�}�k�F	6Rq��Q�8���J����~��O6��� �~EF螸��>�D��+�吐AeTq0��FX��
5g>֞b��i�f�ii�5�II�E����.����9]��&�0�;���(�G�oB.���C��\�+z��w�tL�G雧%?w��}�7�E�n��Z�fc�������CQ<b�Źs��5�;Q���)���-��J68�O�]�f�E.�U�ᛣa�a�}����R��\��I��YS�U��߆��ޔ�U �䴒2�\���VٟQ���
����Bl&��Il�w�݅
���JI����}O�O�jQ��G�%������=g��~�JpRA�L�i3�N�M,U�Q��/�\�ov�t�hfS�C,�����[%�TnUE���p�u�m�O.��s�]Y^�ڼZg�)����V�>I�]�7G4�F��P�����A��oÆ�p�����C;�.���T��x�|I��ν6p4pA` �>8`�m����!�.�,ՊE��9<�� �Q�M ��\�I�W�q�$}��;n/��	�"�|�e��2c/�CYo�����uN�,TO[�^\�S�\�}E
�u\%���^�.ª�M껨�Φ_.�*jF�P��/� ���C����$W�N����YH���>�\Kc��a�V;5���\�5��0�����X����������chj��E�6�N܋ E���Wp<��%�K8�3]��OKr�M�g��T�����"FK�w���Iqmsu���n�8�\Qš�-<b7ƃ`�K`�̙����Z�Z=�����U��u�F� Θ�#b}�KLY��±�/J�nH�և��}��[&�w�+G:q�%-j��B�	.�1_����6U��s�}X��ϟ��ș�Z�������sm��#�J��iH�֖2�4�<ɫ��ˋT��ZG�PӆO�����A�t�:����� R��s�}�(�z��<ϗ� �y���%��@�7=��6$&�B�^C�2���������mJ��yLb�DQ��|���5r�?5��VT��}ec�)��,
�S��Q3?W?���͘��Ӕ�Ǌ�Fj�𲡋��l�����)r���b������5M��o����z��7H��ٝ:�AB�C���a���g��O��N��~����pY--��~K��G V�<4�j���7g�F�eZ�,z�� .��:\\�g����P���X�Gi�1^ЍƗW�L�������:P��]��!���2�����ȡ�<��=o�������5G��ҁ� �
y{�~��ҿ@讥����#,q��Q���4_T�!j�G:f[�/{�)��v�}Dc��1
G�����w�_�;����j
VB�5��HT�Q��1����^,-t4}���=�^�i'Xly[���ף�S�:��^P��������i��Tv g#ⅢNq��N�x�{n�!�d�;��?�c_��3��(�Vޅ�}ӊ�]I� }��M����`�+��2F1U�#Ԓ��5]M���~iE�K�p�J��<y1&<<q���!����O*\~n<3��~n-�m�3�,k�@�e���8��%�B�n���8��p���an�V��d�pš��c����q6q�4��	}��,殺�-�)�/�� ������߅�מ�M]��n7���W �i�4�:��RB�q�lK�·�Sb�}*�n]�Ib��0T輁a=[L9����h��fF�o��5���۾$L�=���S��<g��ؿ|W
1��΀3�%0�F�������G��V6:R]�w��\r��޿$����_���
3�A?&��EQ5�����>օt��ofF(�;؊�JԞ׊�sS[y�/���ˡ[�x`�~j�7T8xB�\���C��잜�0w�t�`��p7�]��*��O���&��O�u0�\7������PY��B�r>푁Q{}c7wA�.�4��!�������y����j+�h�۟x�s��|t�;+9pxc�,��T���� ���\�m�	��G8~'@2f���F�A^���4}�{���m�X�L\)��l�S�k־|
b~{;���/�c]8i�4���-�/�<�9��W���~A\X��ߎ�}��������6}�uzz��I>
em�L|�w'7P��;U�EV�-|�m��?`��A%��v����I�?H\`h��o�{�ݔ�V������{��|9�2���_�l�ՌT/g�-��6�o0@njC������F�`��No�kSU �������P�,���l�%jG,��[+����RkĒ,ga���!�������1���z�Kd�� �i��#�vS��P(������}N����Z |!�E��\���SI�k��|���?�)>H�4�"q�>/\����(��9(rthw�p��%Ay��y�W���ny?��&p(������+�׍�1�Ν�!Uf���g<R�h��	v����<"&M���?31�{��~I;�}�ѡ⧨��Kr�6I�0��q/����2�d�[]1YY��3�؁]ZDP�d~�6Ū�hN)K'�a[����
����V	��3n�JouTo�$::����N����5L'r��-�`�ڝsm:@ld��h�{I�"vJ?Z���m�DT�.,?
���_���/`�씦���o���, f�gg�y7���SF�j���*�l�r�66Phyf��5���<���@ø%�h�u~p���z�f�4P��?�c7X�e�|��CVw��G��O���+�y�?WȾޔ�]]��f��� ���F
0�1���z�:-j�����S�~�U�҆��/劃{� ֖X[�Lc�<�jb�s��FH��̿�/5�?��( Z��p��4���-���L�o��� ��"�?-Q�(y�����{�NXcunc��8������b�t��D
BHY'�PJ����߫9!k �m�Ԝs�%�q_�Wm*\�o�i'���7���
1��Loi��-M�����Z�t�Ȯ�2%t�J_ �%kذ���΋���G�.7��S�FV�\�`��׺�R��qM	�zI�қ���~�Mu\��~K&)Z�m�,-ψB�Ґ��R��_s�%���v���_�c�wX���q�i|J�r3�~f����D�r����l3	<�}�]u]MZV��h�����?�>#2��n)���$����5���į�{ye8�:/̳�3���t��ܻ�(�.T4�>2,�$�6�ͬ�w�#ߔ4��Υ���z���d������>�]��_s�3��� ��(Y}kJb�]�ߪ��N���L8���U�d�K��q^+�C7v�=\����^+l�X(n:�Ͷfw���+C3��\���]���߸,`������,Ҋ�!��WQ��B���G��c��=���Ш���ŷO.'/c�J7��Ԭ�������j��ԭ��R5m7A�>�@��M9����цjk]���N���W*aP��% S� �Nx ;�G�gw>�>����y�p{[�!���!��ပ�WOz,�(�T;
���vv���dI�V&"q9�86Um�թ�9�ϣ�O��y��j�R�w�A����_�w`�a��:���g�� �s�nx6����9���jF��l`�_)��
���\>�ߠݯzu���+
���=��j=��8jg@�Z�ۀ1��;����f=xD�CV�G��R}�1��oK����A^�ܷݔ������5f�f�~n(�`�kT�3ս�4l���vR�sX��/�i����<����Ԁ{����	6/�o�����2���,�țwhM�?��<�,�}��=�*�B�Nds����È��5� ?�N�l��ǑO���)l@1���/@�>/�E5��+�Q�ʬP]XO^��?�#�V�d���Ke��:�,@`�0b~Iخ7�[UrA{d~/Z�㋟��s�	�%��
�0� ���S���x;�����_��$���{&���r�|������z@�����^ؔ�{T�Ko���ʦ7�`�{{�}ox��ϡ��=�0�|���2�z��9�;q�_C��.��HZ�RU�X�v�IgU�؉_��	��i��������+=�?���Ud/΁G<�F�6��FJ�-��WR����?\�<�:A׷���6{�I��h��nOߺ�y�9�N�k��uv0����-C��^�2NXy���P�ls~�r���Oxx3���^p�����cl�d��<ĬeH|�V��0���=��	yX���!v�p*[]<��u(�=�����u�'p��%�o�Xko�q~N4����oI�)�u��>o�����w��7/$毓j����!5-�+hP9�8���<�� 	�<����@�Ojy!��գ�Z�Fվ�ZZ{��0��]��YH�L4�K�+����)k�o9��Ԛ�h�;b	Ɏ9X��;8/4~5�����i����&�`9C��������YW>ffda�M���V�7I�`1�H	�x��	c��� �!����	��?g�֮.��h����h�,��z��{&�͌/8	�y:]�3W�`��GwR��)gؼ��:�b���GdG6�$��1u��jR�7�-�X� �rk�iŀo�kt Ӳ@��OS�-~Ҥ����rZ�2�]w�f^@�E�!�^q@@>��}.�It����ԝPT������@�M��/K�V�2J��s݇=�cN|�́t�7]�U��n���:��إ�}�rn����0�qm����=@�i���z�QV�� ,�i���R��r�d"�8J�*�x�.sDR�hŤ�a��;8x\�'���8��>wWm�Dy�R�&��|c?!�,�Mn������E�ض�`����b�-L�
uq�z����g��)a3���UZ�=(x�g-���u�x�)n��D�I2���}�4�[������y�?�ȋC�>\
C��g8����,W
>�t� ݩϬ���~2@�<�&vX�Tf�^��N�`�@�d�
$[�����s�X� ��;v�=�s^�#�+$��G��\�U@M[�B��1��� ƅL���&�%ʐ�g���d��c�o��P�2;k��'8�G�+���]��T��)��n9��ڐ����[3Q��,����0l*\Adb����h���5��[N��|��SC!�8���V�/��Xx�����'ކ��/�U�2'���2����~��AeL�R���/��}վ2�����@!��z�૩���9P.��j�#���*��������j��lۍ'�Ȟ^���ʃ������d5ۅ�/��̦mg�+:��~�y�S|��=*.�FM묖����,��!��������M�Z�唭�ޱ��g�J�~eۅ��̥x`R�J̡����:%��s��1w��؅p�e�}[����p��{���@MM���D_cM����#�$�M%��ʲo�m�L�uA0p��m������c|7��<�\���r򞩮]�b��$6��ۢ
�����ZuSqzr�Y��	�A��W{K ����լ���sx�1 z�ǫ�������I!��7�/0�*�ت��mguϻ8[}K�L����O
�<ɟ��I�n�aU.�s�$����m�z���ک�����:�q_J��̗��8�����<�?l��g�a6��Wj	��7�'���z�謵�V܅��>�;��n�Ĕ�����{e�$��c�K'((�ɢ������m�*�և�c�2G8�}:���H2-�H���.nj����ܙ��Ofo�]Z�b {�[Jr͓sjK��"��׮�O|#bE����e���]���]�=���B�	�0��$�J����Y�����̙�j�c�X�aN��yX�=�A�p0��z:O&�mr�z�]��kewi����-z�Y�=绹1g\l�v1��*U�J*��d~r��\�����]��|J�Ne%�k3-�T����t?�և��-�˙�1m�u(4.�C���f!IQ�4�N���~;H���no�0�/f�l�t�n*d!W���OR��eYq15�~~]��V{��y�,�Wȷ����6��w���=|h���V��B��Q�D��[�c���$m�*(���i���5tG��ť'퇻���b�\�:ۥ��$�$���>���]l�R� C���P�#;zf�`j�@�K�J����$v(P�Ӥ�ec��M�X�,�}X�)@���V��*�����}���<���I�K�QUxj���=b1 �R܇>RO�������	~$�"�=o�CT���F����� �����}�������n� �U�� ����4P��<�H�C��|J�E��z��;��dq�Q'�P>�a�q����&b���ߺ��m�>� �T��r�YZ7�_��c���ɀesaiKX*�Z�2�W��\<X�K�|�[5��hA�kHp�4Λ[�ٙ\����K�~4>w�Uv�^��0�Գ'�X��c�p��GA��H5���G��ځ&�h�s^�\�G�1m!� Q��j�u�%u�f���yi��H�EV�~h�q�8X����X�؈�fpH��u-�|5��+���nP(T�T[y�cxqG����ωS�^-W4FJpc7�9�1�����xu��Ǌҙ6��G�p�T�a���9X�W{���$����vo�zs�zx����)P a�έAC���+�@b��F�i����y��w 2��K��z�D� =WE@l���#���4pe���
�P$% �F ����;��p�e��ʓ6��;V"{;1W0����$&Fzk��Ĭ���o<���e�`�򱂑�:��&�p}[/��Sbsn�4�u̐���EFH5Q"T�N؅���3�?�Qcl���A'Xt��H��$kV��"U�G����W���ݼ{v`�R8(lŭ3��%c$��eH�P��x�`{��λ|�H3MJ�=�~�.\t����R�e4�4��e
1T=�����i�B�[�E���e:�1��H�ȟ����Lq�upR�-!�<x޻��x�����U�w�<`Y�����!5�vCx+.�I�_�����̈� � ~ǭ��ndg��^EV8�͘V�T�~���)<Pq��p1���c�|qO��A�?�A����[�ŭ��T��Y���I���K5ȴ7�_��C'6��^ޘj	�Ul��[S�T0&h�=�U���0?��,[�6�/��H����1��/N%��s+�~Ni�W������X��7�U���Ej~oZ�P��Ф��,��b#�(�q� �s���ã+32��>��قe�Q�į{����w�ݑ�o��#'Z.��~��Jh�R��̓:yӫ_�4u�ټHÕ�e�MU�'ͼMR�Ԓ�0�rGT֧ߺ���1�K�-�R�ܼP����.�F�ĭEZԱ�[�ל����q�W���}�OY�Y�H�6�I.�>���#}_+!��^�W��E�qq����L>V��_<"��J���?w������+�x��i}�sP�i<�'ȟ����������.9���iC�>"��[�ދZ��X\�+���?���0:�#@I��;�f�X�Ԯ�a�r&Nkɷ��F�D{Ֆ�na�ar�WP�X,�JT�顰�Y�) ;�8�crz�H�J������y������XHQ������20�1&�3��v��H�Ģ���O��@ 䧀Tqة}+�բ�3ϖ�ze� Ӗ*i�/��e���c/I�)Vg�&��L���Rvj"�� 0�Ƚ =Ǚh�����V��jP�QWY�	3��Ϛ]Z�g�����;ws^B�)J�gʕ�v�К�{���u�',h=Gm�״bG�RY2�+�]p�3eGg�J����}|��7m���gGͧ���ڝK�ؙ�o�%�
���fI 3��9�P�p�� 5�9a�T�����%�߭�~����y��Ì
j�e����zo������xN��tU�!���	z�B"���z�䴖��DX��>=�I�����s��02����ٿƁ:�����#da�ջ��S׻	o�,_!���j}z4)i 4�<��>Rei��2	F9���L����)m3&�=��vsP=9�]���d�\�6pO�L�g*aݿ�J�&�J?����D�x��Z��d��Y�b#q��
�L�������54��uv�^jSjb5�)!�*8u����de�M��L�痊NQ��8�T��J0*>t�����;y����Y�RF��&&���������{S3C�7	��N�}Փ Cl����!�w������D��⭣s����w?�vŨ�p����_����=ѯqEANh��p�˘I�`Ԃt����Q�{�};���A/��5�eTBc�Ă�qk;T#'T+��ƶ����m��9١Jz��r�$�#��ܵ�ǎ��׸�?E���q^�j���,q���Y�?��c������@�P��i�vTݯ����]"�����R{���Hɒ0�y|2s���y3�TЩ����9�g�2�s�.1�?U!���o� �)S��9�GD��`Ǧ��Rgu�wl��ρ��-(�mw�����)��DP~J����h�c�3�U�L�{Փ�nhTK�q�K,��2˫Q��������c� p�[BŌ�o�D����%3Gʼ��Y˷�Fo�K� H�ޭ{�#4���D�vz���ըa���|ٜ��(�����JbC`ay��rL��(GB�>H�c�� �SV��U�R�
���ß'�Y<{����΀O���6&׻��Ӆ�Qbnb��w���,Nƅ98G����5��T� _?Y�9�qM��oٰ��R0W��VW7� H���RA�����o�S�~�Ο����g��x�^KY�����N��0�~h/����0¼�ْw���=����|uD�>�Ⴖ2T�&pQ�HJ�dt�T���)<e��b1V��u_8� A%�R�V�?��,~�v�#�pe<���Oʺ���/{�}}1�9���u��ֶbBf���3Y���bK#g�"�s�k4��o^�A� ���&�>:�=�	��U&X�����5c*�Veb�`	�Hڼ�K�n��@��|D��+�똑���������Zyy�t,�*U��p%���p?X�"?�(�?`M�A�~h�#���E�?X��LJ�MI��Jг|���JeA���Fb��|����6*�DNefż ^Y[ՁGc
��`��KV���,91�E0@0�]Æ�R�MU�H�|@��Eo��$��~g��}sp3�XY���kE��t�%o��	x4=�Z\�h����@���S�XK��^5���2j*Ɍ����С��_����B��!��J��D�n���@u!���Nּ9z|>���&M�u����0-}�����z���p�&��Z�P����*Լog��s��e6�\�����H]�CX�~�.��L����ȼ�g�n2�ﻖ�Qnh�Ժt&�.�qh5@ �_���Q4�����3Q�O��1�
����p#f㏹��\4��Tc%�0F�>�%�\�)YI��q�^[L��5�EG��֎���C�w�(��;Kl�����ɖ鷛�qo"����v
J�C���F.y?QB�X�^؎��:ή[`h����<4x�P�Φ�<&&�yI�[S��/aJo��OiE�QTb�L\V��{rG��|�����9�� �	4����vCW�J��,1�}�JUp{q�7�M�%�u��Ҏj��L���=�B��(���z9�y��{C�9�j)D�=��/m�F�G���/�;�x<����&���Į�I���lbQ�0�r�*Wŝ��<�\0��VX��Q��g9Ce�-
ì
m����T˄���FC����EZY@�����;+/�y(��N��&�&3d�8?�2�ȅ*�_��%�'N�	B4�|)� Ii��
;j��,��̨��}:�08��ܙޟ�7�G)��`jMll��'�[;��C�S&3U�;��n\��2�G�8+<����b>���4�j{�	�"�݊��37oٖ'j�C���^o�)���nb�Q���2(�����U6�W��e��i��89qF��I�5�E���.��P/=�P��Ul�x�J��t���hD�X�EN���>�ș���\�WXۇk�~:�{Zc����tC9c������K��5���N�C� �(:P8A���(�R~��	6��Oy!-�3�(����9#dB�F�D�v�s�`��A�Ml��VX�'~��F
N�D��M�����J�v��ES���/��z���EmpnмP��O�Xm/X��jd���MFKgv+Οiڛ�^K�N{\EӉ�*;5N��Ti_�d�
�E���ݜ�Z��>�\��=uP�Կ���f5�,<�K��q(���9�W��8'�*���{N;�>�wb��>�m�ρW�X�4�j��/��i�ݽ�$�V�k�j}�oʞ��n��WM�+��m�.M����V����@��4a�@�fv��6	���0��*��/�|��z��3���YCP�@h���]�cyd?�����;E��rA��3�E��1p���s�����G����� �'�L� ���j ����0�}�x�O��`I�����a�ʿw��B@�U�`�;��ԃL̘�z�����OT�d��%>2Y�m�>ۏ��h*"f\�����x�����5�GH�aS<��{˽��Qd�H[Ţj��OW	vU��������5z�o=&���:`�*�}5z���Z
삥r0W�0�l�D�I�*}�ueT��4��[mI;�	����Uʲ� �FT�(�a�G�iS+��_���! �Z��� )J�)�%?*
ީa��cX�D0��G��r��f��r�*x�&}�>��`ٺ(m��R����}8�`�O�`\��dSLn������pY�]9Q,P9�g�
��~Sy�ls�y����p؋�Ŏn� ���FhC�F$��433��cx|4���YY"��jq�L� 0��a?� _�V�>p���v��݋lv���d2/�����юq���Kb�a��>KܸƆ@-����~RZ����?��&x:I��F��5�^��ES<�|����Үt�:%������
�@�dEY��G���ܜ�]�U�k�p2�k���02��Srk�릢��!|��mYz ���M���Z>Y�jMd���2���L@-O5l|,?�P�G09HB���^�fب���ax�(ٌ�����Ոb��2I�G��ӨƉ��Y�ԁP~���e_Oz2��Ѐ����^�h���ˊ����Q�7jj�h'8C�7�h�������̼l�����٨�7��_�r]O|ǉw�w�*o�s����ߣ���3�4G�Ź��p[��?��g=��%i��Ě0��y����F��
&h=��`����g9��[P�����2N�Rn�	*�ʙ��f��	,F)�a>�XUg4[��PJշ���FY�qvX >#&VS����k��T�<�N�!��ɂ�y.�ubO6�P%:�A)&6���]y��. �}��q<��R�o-E���F���ҟ�>�F���<8|�7 7:9���o�ǰz�,W�ѹ�>k&mQe\J�ѝ��D�ЈcC���6TeL�'g�}[�(\	s�c��"Ȝ�����Uڒ�`��c�y��ʂ{r[t˥̾��&c` �VIL�x���Fh�������2�:m���q�N��R�Ȍ�^B5�1��E�G�~��&}�3��}����Wțe>�V�]��A�/���ˊT}R�J2Z�o��c����[SÏ�b=���=�
�~��}�,�z��f����i�CbnSw���S�������)�e���a��NZ�K�ϤI�E�ĉ�O�)�؊�2��� �xo&��Hހ�:�2���z�غD�lN�m���:,���l�2#R�C�eS�`�����WLJ�d]᫵[U��4i�����QQeY�p9N��"H�-((ݠ`�
J��A��`���%��((��
P�@@�H����
I%�P�(�=�ܺ83��������Y�캧�N�~�ާnյI8��!�A��J����"��~R1I�솜�w�|�b!�����L�D�t���z�L.=YW�3�|����q�O�B͚o{��J����y7ﲛeV��V�1��p�g���]�\[�u��l��jƝ��ؐ�"��>;��R��sb%P{;���6:@�D�>�*|v���Ws����|9�S�fBMz�
g͎������Ǐw����M�FȯKm}���ۙ����b<���[K�e~�l�@��MZ�[�R�B�`]�j�Ǩ�&���aA��5U����"�@o\r���'���|ˋ,_�9�/F@C'�:S��uG�������1�LT���/��б*���NN+�Ӛ��W/"b"L� �aP��Z*��ƀϘ�D��K��1>����m���_�o\��`�ᣩ��"Y��x5� ؄���j7��|��~R���rF�l���`�rwJٛu�)%�W�|fS��e긠M?R���+)\lST��v����xh��.�K��:�s�B'�x�����LVS�cL��|�#	�e�
��WfWz��ښ��di�}�Xaz��˸�AT�X����<\����xY@Y����.����+���f4��Dwd9{�����a����m���<��B�󄴧�gظ��+�/o���MԢs1����R�
�t��v�x��naU(�'#"9�3�=~u"����}#��CQ�C򩣔��"фn��ya_�Q�2�Ⴡ���"�!��:��z����+g롻��vY�J>���9[#$���}rB��}�E�n�F7&�;��+�<u�p�3t��z����%#���j�g�q�R�p�ͳ!�����k�/s��w5���n�io�'z���6���������5fg�К��慬�Z�{҅�4w���/��)�>n�D&�����kG^֏��,����poI�����M�v�?XM�r?��:����4j���jw3�m�m�qeN��zy�4F���U�"0?(���	�s�v<��,l�q 1�)HQ'ݬt}V�t�8�`Ej�_���	�yq�
Œ��= T������4<ߔ�E>+�e��5h:��j���."ty�k���{�qrs���'ݭ<]������0�),����gh�Qn��"
���zw�m��R[���F���*v��8��k������Gr^�D�ls
Wy��y��^Qp�cX�5h�c}�����p���u�����Y��;��9P(�/�)w*�G��1�'���f�H����8�kj��(���i��*�ӏ[z�DLz#4e#��S���@��Ͼ����:]c�Zg�h�0׾D�"�h��z��W��w���R4UN�)�1��i#���Ҁ������CEe��NJ;�0��A�6��E��zW>�\��Z�#mU�&�k��̳�v�fҳ��0^�p�q��lKp��9:���,ȭ8OH#Fπ��U�<㧥��a��S�^yu�F9�2���u�;��F�һۣ� �$6���������͍mor|�{�P�c��3��S��x�b.uc��~-�iq�]�Bd���]�����ՀJT�꼀���pM��pi�'�+/fl��}��l���� ���Qv��-�j�Y�(F�6x�Dz���!�	\��n[�ݓ�%�q=�B��Ḟa��_ ��nμ+^.7[����W�u?��c
�b���c%astPv�7�e��5UgT���'�����,�G���^�ͯϳ?}/�W�B	u�ݸ��M�~2�"�3���]�����	�>�+���sz~�*��2���+����1}:�N�䩛��YgX�̌�`�u�˼@&�{g?�0�����:7��A�Z���bwa2�E�B�ʂj������\��
�a�B�cF������=��=ν��Eh-�ܞ]��M8��t>h��ʼ�њ<��;>�|�X�T�f���h������`��~��צ�L��.�9my��5�'�֠����E�<k\(q�h������w��Jc��_`n��Z�)5['�>���¼�lwƳ�Z��2u����Y�~��1��=�S�ݒQ6�Q�{�0׵=�\'� �[�r<��-�F�5�o��f˟_|%P*���#O�P#����HѴ�ò�����wҰst�W�w�0�E�(�y�W��%�U?����J�Z�]��˅�.wݰ݋������)*�Z,M.|�����m�]��ȓV���*�!%�n
�
���s�P�HF�9>lwxc!�:,�v�}8{{q�FżZ��F��,� ?�L0�ȵ�҇���G�%N��8C���M]�Y�����\qo���8�r�u:���4����X���.�"�6 ���'΢-�����`�T�A M�~�z�U4o)U9���CP�$��3*Sx��YO6Ep����.���7�j�y:��U�+ZT��gTs��|	R�NNЉ�Ivr�є�ީ�4F���eV
�����C�
�%���u��z=^H����C�����Nkj�
����f��aa�g��`�܉�k��:Hq��5�mϰ���	��ڱ�	����!�X� ��:�x��@���ʹn�u4]l	r�xz���o�g��%cx;���.�(�NG�F@��������4�I��tIy�hW��`[>#l��@P#t��&;Y�
j�k�9ۍ��������Zt��`���k����:�D���m:Ʉ�*��̲7�d�6On�P����#T8`�L�j�P�V(�]�#��;�g��aq�SQ���7q;�I�����q\ͭ�Z�~`X>$���6!�m=5�_�2%u����znW����@��e����Z�_K����%�sD��Mn`5NF���I�*v�O���t����)O�z�η�/c�������8����5�������X��-�쇍i���u��M�8%��Ɋ������s<�Π��p�} �,� ��mU�Zâ�  5���6�V�5��("0nElJ���(b꾾�_[��Z���;�ɢR?�C`͡p�SC�92�&:N�D�Z)�,2�AL�b�k��Y0��4a����g�ݐ�5��o-$)�^�GjB�e��Nmw���%�-��IX�.�DL(e�~�����s
>d��&�m9�RpFG�ܼ���|'�iv�Q�B_��C��L�N�_OS�-p�zd������P��`{`�s1�4�9�Qǎ��Ԑ�t�#��c�GF�g'���gG�u��}�<���]^b�=�3��{�����[XwGYz��b/=���I/�t�䡝�"��L}���%i�ߔ}�����Pxw�}��^X����'��E-&C
Ղ5�܅�����dY���.������ݗ��^�oـi!�����Ӗ��\r�;��!.�0����f��|"h�k�����h����\��,s���:��n/vʱ<�k��X\c^6s�m�9��������sH¾��7<,~/�M�� B�ܘ;3�$~�z�M��?l�����;z@ӑ3J�l];Th�>xC#a��g�9�[`k�kZ�<ǹ�N+��}j����k��[���=�,�ry\}p���H���(c���Jx��y<d�wa��I��ɸC��]��Z��o+�ο4�y��d�<�Z{���t<�Nmi'�c	��GU]2�I��Ȥ�����}:�����sA�Ōk��W��Ż�"_|n�����X�6Ӻ�e)�*�
����^2a[�8�P�$E�kh͞}r��Ǚ|qqw��8�ӑ��oP�qz�u�&m�]��-�Ƙ����"��7���R�I�5���y�ft��ΡО���,v?�9Ğ����.�q:��1x�Ξ�/+�1�$@���}����ڧ�B8Xٱ��1�����A���z�`�t��}`�&����84zMa���p�h!�����@9^q��Y2���V���}�@��'4f��>o���@����^��#x2_�AN���RT�e�^4��7a�]i��i�C�{Dx2�|������U��z���	�N��,�N�4��	�:��9Y�umo�ƪ>�w?��	�v�}{j��1Z�!��ׯI�~��P�C��^
z9�|���������)�e.!J�i�)�G�ŉ�X �7* ��a֪ajA������U�<�џZ�߃�a���J�w���/�Ã���5��NKr�Y��>��]���AKz��W'+�Ѻ+;�����c�b��@�~��k�1q�(�|P���1b��'Z�k�:V�;�6������.7� �T.�\4Q"����	�)��J�� ���j��\����]Rh���KĜV���Q=۞�uKiK����D����`��B�=�$Y6�:�)���c>�s$*, ���@����C�[�kc9���3�zP?� ����>IX�Wj?{?3|�n���ʶ���I�D�����e�ƿ�����5
�u�t�;��Y8B�q��Z@;��_n�M�l�B;iHϛ6�g۫� �������S??�����Hf~������\G=���ю�b�)�耲�E_���?��d}i.o0~��C<�̀���s9�/�-����-��K�u��*(>ة�?���k�nv�@�ځ0��u7��p�F[n`������k�_ƃ^k{4.?o-������@����6�1um*�˫�_�M̹Г	S�؎<z��3���r�Z�5�·DLt�DT�꥟c^�i�=m)�"����>0���J,̕�a�+;�ڇ�k%5��M��( S2�����]b��.8����iv�+?�~��NKI���[��}�|-��P~���=������S=y�o�����<F;i!�����n���$dk�u�3w$x�/��Gئ�8��U%����؝f��������h A#2a�O�O�,����=my�����B���M�g�-�?��#-��F�fꎃ�9��3�𖻔=���1+��A8ᑠU7�(���=f��Vg��K2Js�;
>����:��EO����`�fm�vD�t���u��a����x+�iԎ�9)����՛ﻔ�n��0i\7=�$r� ��x8]��v�l�ů���DHw�c�Q*�VW�Xd�1h��s.�(8~�0�ԯM(�tK�Hn&�\Je�_̸�8v3/X��i�_V'ҫ���&	Y����6��ՎNWqe�:-[Kr��lC���#���U�;�:��\g6r���]�,��IX4Z�w�����3�g������Ŀ��{^�.����"�*����!�V�����ڜ��9�%����+�C��xv&�H������yq��\�e��n_�=���]+��6ފn��$k�̭��5L��={�����
�����on�O,�ۗ��O�,֍����w+����sRC��,T1����Gqe�P��ç��x��7�e�W�s�x𾯚$L�D���W������e":P��0_}t���Kk�c�VT�~%����[|+��*-0@O�2z�D�p����>�\���o^�Y�d��_�xsq����^��?[�Yӳ[���)R�������^����+�EG5�UJ�@O��@\]]�^�f�$'g�"��(���D��F���
��7'2c���O�N��{���+���y�����|&	o:��Gχ"6%h���7��]�ǁI���t�ʸ�s0���;�|]�eT]h�h���;0���|i���쎱��r��ݾ6[�������מ���ү��k��7?ؙ�^�zc��Μ���"��:�9V����M������کo�rq��f7븓��եz���~�����dwXk���èSB�)l�h9��a�3Jc�r
7���;�o��w�8������%�z���+{�'���C꩏/���$ǫ�����\+�} �x}:�n��i�?R����������È�=ն�J���ӣ~��Y�+�_��Ƹ�U_;`���.�Jѽ&���n5��U�Gf�,^��L0�5�
��)p]��1A%�+!���k�Y�����7�-�;-���Łm&����LwJC��[#[v����h�R@��߉���R�_��k��u(1�����m�Qe�A`�Wz��1!��U�o�?ޯk�dXx"t��wA�dc9}�A�{�S����@>��*��tDS��b��<e�ɇ�H�]�}[b����8^��op=��4�= �?�9[�b�W��e@�7j�	_,1���K&�9�J�n>�.��<������Q�m
emIl�\7�%�x���f���m�r���͋�*�\��jsk�4������Ot�V5�1,�;��o��x`�-$�/�Ә�F�P��b�7���&�e�%�ŧ>F1�J��,:w�<�O3�� �y�1YQޛ�T������݃�=ѡ���h��f���m�
���M��Z��G�D�ǻ�|W:���{<e`�o��֬��5Y�Mi�/�pe�oc|}}a�N�{��
w9�͢~�+��D|lՄ�hq����G�3�����vsxh=yS�{:�#!��^����vB��E�(����9�R%�����J&��zeG�{�E4+v�Z����;�W�9�>dg�4�˿��9Y��q��l|�N��A�����O*�_��Ϫ�M�Ay���Ŏ��iQ�Į��JW͐2_��D{��{������M�T`f��C��[�S��(���|�Z�r_l,�`�e��53��#W��ROR-���[�Jl<J!���7wl�p�/�n�{5���(�^>����!ioNJD�餢`E���2�՟l�3TD�>Jf��Z�8�#�R��5�4�����0�����'���i�����_���)M�l)������!�j6nes��s=Z��+�3���ٗg�Y�IP�/�y��ce��q���si�������d��RQWN���nU��]�e����¦�����	�����	
[P0���L[�~��	z�����������%wFR�,��Fʍ���O�Άv;1�<A����!=�ۂ�R�I�V�/$�RM��0�Z��^��a��?s�T�K�I�VL�ӑƮ�lf�/B�->�l�/��O�'وN�S�O��Z�N�tS��@��rK�IԣV#fN�L}�$�Q�o��8���yO;]s{�cE�y�X���Rp���rM:���]�n٧f���kb�_�pS�<����j�P~�;e`�3�5�r���V�|/`zG����ϾA=7?�()Y���{��.���[��ݯ���Ӿͫ�I����ܠ�F*���Ƈ&n/�L������Y��Φ�Vz฿�˂����b�b���F9�0��}��5�������Q
c��R�%��E��=��/�t�[�Z��z&L�μ��,�m�ut�>��K�E�9u5=�2C��Ç������Ǆ����
����?d��"�)���o}�_������Zh�������������D>����o"���&��o"���&��o"���&��o"���Md�F����W���[���(s�ƫ��n��s֫l��>�� �rY'�����Đ�z?����IOl�����e���������V����_��&��o�	�&��o�	�&��o�	�*��������o�	�&��c�jW.G|��W'����v�v�&�@�����v
�%�K�(E_&����wyU��k�\m���������(ܾ��8�형�lL�����MtK���/��p���{����ȣ�ˮ��𳔓�/�Ô��WyC���`F*nn�_TT�O��z��EWp�g���
5��̢���G���#��8���Ƿ���7ӡ,��7�-�`�x�~��JB��׷ֽXu���p�C����*'�y˹m��jNӄ�@�Mo%j&7ה�_���[��"A����{�a݆��Ug)�����l��� �ɋ�|imfj�^�ݱ�ɉǺY��}#s��c�˨B����O�XK�Ǻ���U���6�-e��?^�&���h%��o��{QRRr#sS���u3.�k�5q\�Y<��ʲ�X��򔢬ۺ��Q���la~ў0��y�����\�Ù�}��e�w�<�j���gT���	�臢R{�FW�zH�����k~OϾ��w؝�[��X\r����A:䑳�w�)E	K[�>������3�ܧ<��}�@�E"�E��[�X�r���M�w#�Z��N����ػ��3,:� n�8F�f�LK0���$i�F�E9!�c(~�'�W��Kz�hg3�;A�s+k�!!h�ٯۈs�����ϫs���^�(��_7ISeŻi��گ����E՛�	3�.cJ�Xl�?]���DO�@
�9��Η'�eD�1�̾�(�b�������O1�)>-���\|~��(#���8����twKKKg�G�&�~4�\�H��m�Ǧ�{�ĸOHJ.f}Fˤ6��:H�?u��f��f�J��+!�O�����O~�Zز�6��HW,�ʚ2z�6�a��[�����&d���ę\����u R^�7���F���|���+�F����{�5^wY{3(NƁ���w#ΩUUUB�h�)�mX�R�M��_�˾D*4���>����rXU&.d�!(����ۜ%:k��)�*�*G-*C�5mڇ�/N����us̲p�������\]��G��'H]�h\��?e	{��җ\TUUW��AW#��]wumy�/%�t��)؂N-�NY �7w1R<�-�as���D��//�uY�L�Ѽ���T�f��Xu���ER�-w��/OY5M�y��`J��������n�Ͷ�3�e�D�d߂��r�5�S��U[UWW����}�e�y{����u�Dt�����3��Oi;1��%L�������^g�����(`E����`�؛7��m[����i�Y� �#q��Ν;o����A�,��&ƽjR��7�2qm�Z���R'qO�o�������gm� �<�������ϕ+�x0����Z$xq�D#yv95U$ ��[h�O`�WF��Ow�1��p��v��+�:�(�>k�ak�o�3v�8�lp�Ό�rqq�+`��􋰰p�9�.�9�ͷ���=O���n�ދ,z��{���CZ��Ζ����i�q��(+�۳���ʒ������G�1\*�cA'qϽ��=v�#D�T��l`�-{�i�����(����9�G�OJJ2�%�`�Nā�K�L��^���S�|���5�
ПgQU�YN3���}E�Q~ ��(m� 0�9�gb,��n�̒u��]\ḇ��;<&��&ɔm��b$�+J�� �^b�oꞚ��M� �	Fh��W�2'ǣ�#�/�q�)�.fx;��wqD�j�@�m%=� �̯�l�Ǭ]˲^���ƽ�T�VgM��~�yA��=afVzw�����(��e����A��S%y6����O�摈U߹�����D�k������OM��n`���j�U�B'�Kw�l�Nn�I_�x��Һ>H4�*��bۊ�"�2���6�@�:��$�+y7pI��`�k�vQ��.2Y�,�@	Ϸf�c ~9��ɝ�*����#(K"���>�\�돸hPL���C�y6	{P�v��+��ńF��Q�p4R����b�A俬6�/�N�k���A�#�L��VWW��X~0����)tҵ8������L`�L���@��������+�z��'�V/���U�� ﹐BٍT��U	���~A�H"�ވf՘�|i�/S	��0��[i���qUn�ḪaN"D�b�(�Z��"��Y䭱�,��=�� )W��4�.k㘪ś��I� ��x��/��ܹ�d�f\Ov�S��aPf�Å4d0g��Q������k��=�Î�Siii�ǿ�,���?��p�"��	�����}f�fà�,�:�=�o!�}*c��L�g���`���S�#)
�q���x�eӭp�"��}�36i	kU��q�0hmm��I��Z��&�y�0 �����)�����LY�(I6�	h���q�g���VlD�3ov.l� t���R�:�[�)��'Ѧ��"k������d��oġ�$�2b�¶i"�򼔔�s�t���]�Q�%�g]���\aQ|���e��I��&G��)M6���&?!�؋�<2�U����Xg����̩�Y�p�$�_tH�b�d�u��i��O�8*Y&x�T&L���}~077�m~eM��^'6%EGG���Z��kp��v;6�p8�cjΡ��&�R����=�m��:������+B�����!i/�y�J�s��Lp���Y�����d�yv�h'a."�Kn��)�ri� ���C}#�ə��P��xg";^
 W���/���򜄬R۸]v�DZ |g�j�Μ�8��̿tb�d�t�^�dG�Gi��
rHx�S��N���F�(��t��D=h�5n�]�R��S�����eP�g$N����B�2��^ߍq"�7��,yiF4,(����'�TE�n�F8`�ƅi%%�1{�T\�B��e&�z�S�&���ƛ����� m�Xޞ7>��~��.�Z)�62ȔA�2��od���Y29M�!�Ǚ�ϵ�N0|����ݛ%�w#*�ï6|����H��<v?j_!��,΋FN�_�Ci^x9&*���,��=6�*@��d��U�{Oq��ރG=�n����B���ߣ��ֲti�����i\��W���9�'!���n5K�Q@C	9I,�ȅF�}P)?���㛒zt�=t[��c�TY0��fxBL������ǲ,���z⦪��R���T�����ZSSS�g�Tg�X��g%A�蛙�Q'����mc�P�ؽ�Gi҇�1|>��S�$�wR�J(n<{琢��i���x�2V�^�N�,--�`"� ��+��v��+�A�Ӻ��u1�i�.�zK���5З=���� 4��Mi�� %���{OyA�sD<Sx���e�������kݠ�r@I^a�+4h�V����,7ۄ���j*��[����n�6H�g>�u��k�c���7�>��V��:��|/"�J�.2q�4���x��:;n��s��n�����>�|J��y�֌D�La.�"�'��R�	PǸe8�˝��!�
�7���<�H#	H�l�&
Q�vO|��C��6�.J��q�M�F���""͐�[��"���*�n����y�b�Ni�a?��d|3fX[#���&��F�}T\�#Җ�l$��<�j7���ꃲ'�J"����X�Ƣ9���������I�0��͵�Q���~S7V���2B[(W�Rm���m�"Ng�gC��<��]�`Z��v1O8�d�"k�Z��z�)=�PŮ��w� yh0ªk�gS��֎"`n�����y[�W�3W�͇�)M&��
0���~��,*;��Y������VDZ�\4�-�X|i��Y��r#�~++��$��@a.�Ir��|��r#[�!��{/T��N^��ld�h�}tɑ��7���/q(�����d�x\is0��6��)�K2J@7���ㄫs�LN��nwi��A{/������&&姱�I�^g^����%IԴHI��ӳ�ެ�PfB`=�.�27�,I&�������e���J@q�!�Ҟ��^�*6W���V!�@��-�jծ��(T[M���D�!�X�����m����Y��'0�D����g��FCM4��Q����ޗ�>'���ĺ>wo@�b�ߏ8���+b�M�q]��.��X-�٘4r7�f�	S?�b�-��yb)�s���j3�ld�S/<t� uU��)�%L�x�TD3��<�ǒ�Ⳮ��HW��O�L��.��=�ʍ�Q����§i ��LL|W���_#��<0��/��Ҥ�0 ����n��FEDA|�x���JT����u3��4�2&�����r��h�eh�M�z�%�dܹsg2 [�{��ø��J������+E�X�l�
	�(M���G���6hLU@�.\w���T��S�D�n�V��"KS*��q��W^0�8�F���������J:''��)ER�Z�V����fyJj�N�<<:a$�N�-���1K�3�o�`i�z�s�����m�����*}�6�]id\5>M |:�g�'WR�j���X��aZ�uO�Կ%�(����У��4�NBz�3��\; w�^����9���ݩ3O�\�8b���������%����;�t�@�e��2?>>�?Q'-
����U�8��$��˗�	�'1vbܫ$��$<�S����6�Gp_6��O)�+�gK��gH����0���;���c���&���R��OP:n�}�۵��'����kl�,��
O*v{*�F�\�6n`W����_� �w�2BQC^�������	l�T�x�΅��Ԓ��p0��fC�Ջ��3"�$`�̑Dq|���FǕ�����PR�T#����BZ�to�Q~Ď�dބ�4a�?:�2s ����6�B*Lbx~,N�ӕH��By��D�!�>�vۍ��ٗ�-7I#Ch��3JS��j�6�N�ҷng_����ݒ4�'&I;���ke��㠡&�� Ȃ�巐���@��/��07���F&`T��xc��}��d.,�qw� �Dժ��<����e�!�ۅq�Jh�ܐJ�򇩓�x}�+5e��7�6m�m(���&S�O�c9���8'���A���z/ GO���`!���\x��? ����sƨ�����D�?��W���8����d�Y�
����8��Q m�j��`ⵇh�nnn�K�������^�slhӗj��,�XIM�Xn�V�T��p��:����q���ڬ"����\vƟ�;J�҂���q�6:�y�������>���"���d�/�$J���W�V츭Z�B����Z��\�BT�e`�Mc����(-c>��ێ���I��7��o�\�^�+�ku�!�k{`rr�]|BBB
g�'�3��d�)3k�C���o`�8��J�y�����P�ո/c��_��@@E�L�F�U�/(+��5j�8�|AgK-� Y�4	��á����tn�����:y&�W��IQ��C���n�$��LC�6�+�}&���c���6H�cO@�yaÌ��\8���S�ƦqW���^K��'CCC���rK�_�Y����+=s�҄��<�Vttu'�;v`r3q��ϟ?71�����+��<��Kr
�j�%�s��C��Aǐ����y�$s��!������K	D�j�휩�-��(TX�:�U[�e�@���U�Fh��z�VE��{�@ ؏f�Ct�%[����?֑��A�>��+�(:2�����\��=IM�-�y)�Ҵ��s�$&6Vv7X� J~NR��o�"�2B�/�5�2%%��8�@��q��K���B~�\����%�6�?����b�%��i�0\����h�,������(-q`��o/�Ft?�Q�� yj�B��C[[{�0mN�u�V�f���&�V�[qs�?�z'�I>�m��ӟ0�\�Ч��KN��d�n�ֻ���㜜���$���w;�{�YFT����7���C7h����Nt	y0`�����U'�&o�cw�^Pwʓ)���k�͑�p�8�醟y��P����Cm���@C+]�z��Q���h��k0muK3� ��%���e|+�2����=�Η%%�M`��>a�Ά�m�-���3��@V�`��b���y� �%��2cz>jB��G�`��Aט_GG���R�ص�"���](�W���U�_60X)�4�A��/��f����%��Φ�[���\#%��}���4C��C�|�t;�zz�Z6��쮕f�$���.~<?������I\#�uy8d����h����e`���g^� �=�ow���z�о�y��U}}}:k�d�,� �[���鑰��E>�tL´�r�"�>��.�x���3Z$Q�ç��z�$��iw#.���D;QZ�Q���{腧�(��N���M�6�?ͻk(��ێ�O�C��~�� R��~
&`�*���DE˽mm'������(l|�w�V�$�&�bb����_�;<Y	0[m-)Bk�R0�����gձ���	�1ץ��+�� ����ˎ��z�GH�Gz ����.��\ns_��u��cD���k�-ΟQ=����e1��w�_��4���+���jN�&����n��ݿҷ���Ͽ�#�I�q��gǘ[�6J]��:���o����w��=־�䛜t��@�XI���ť�g�tn�5(\fb�%/��B�0O��0Vx�?CB\�#gv�e�0�(�\|h��VIՌ����(���<�}�����b����p�k��/�����qq~�87VXX��:���}���b���;��J� ��=>�������A��$U�ʇG���g9�ui@��wk�t�l�8D�w�����LΕ��ù�
�+�q�@��5��L Ns�@�$<�ʜ�9��{3U!"����%�e�_'п��1;J���i��Ũ��ַ��h�G���R^�J^�`n�(��.�`$���:=D(��S:�=Ϧ��l�*	B��M~�832*j�"ʚN���ƙ���YaU���2W_r�={��H���v�����I	�`Ȇ'�y�7L�͇����q��>���[�'�tpN�4&2��UN|�����D�Fg��f����5RM!R�A��٦g�f#K�Lvq�������K�ž�v�ymT�6c=�Sj��
�P�jhl,��`�FA��8��\��I���ir&�G�f\ll�����Rt�����4]��T1 �64�bk���qa2�9k�٣��4mR&:巉N�|En�����v����DvQQ�4�z��?����N�R�nL\7�.�u7$<\��ral�)}a����C�t�l��G(M�Q���b㔦�ؤ�V�I�b?�*v0i,P�8T�ґ+i�n?_[[G�#�~C	�P���V&P�vD�E�r"s��Wn��>*�r���K�?�Tys�뎹,�l��W}�Q����Ck��b����r��\_��vS�/�!͕�:=2��~�.���b@ ���N��7S}��=�MH(?¯�����P��EP\���n�5>m���Q���R�"(���x�-�f	�a��7<��c��t+|�$EVΪ�Rg�_�N-w�%hABټi��ߟ�(� m'X�Ej422*����C���eY"x�L�U�d"�8Y\�� jN4J��s(��:i�K�VM�I�Z�nr9/w��Zrs񔕼R �]l��R� �-W1P�ow|`ίk*�	�߅Y/��Tt%��?X�}x��xr+�E���H36:&�H$~�AP��e���yү$����Aۼr��=�h������@j���A��YZZb����� �j^�'�/A_R,�r�1,�.��/�!���� ObX\^/�(����@SX�.��	��ﱵA��\�y����6OT��p$�]��f,F@���lr���7#-۾��)��Հ/�0�ڃ(M� Y&G!�g������u�̍��Eg�9�Х������/^5l�;2q�|�t��,:�ejl���Q[2���9	��" x��;�'$%���L�m`Zy��]�u�K�C<...���U�|�#諹����C��?�X����j����62�}X(W�D��}Q��} ����CU�2�
�Eb�Џ�!y8Ya�@���t0VbC��X[��{J��
�Z�X?��y�6�J_�B���]	u's�t,kG��^J	r����2��2J
-c$�zJW((ӄbYId/�qU�j�w��ƺ
gE����I����ׇG���h�U�Do�FRDDĤ�����s��"E��_'+W� ,�� ���zʁ�`_��҅٪X#m��3[�0XWW��Jj�~WkHjjj�J%��e�9���޼�\��7:�6����V��K3�Wָ�J�\~f$␶���w�f(E$õ< ���D�o4�D�7���Ci�����ح�(ÂG}^|ޫ� ��&ps���U���g=]XX�3�7:�<���y3�G�*��U��+D�]���B���
@�%Q�W���ǰ�E�H�.[�/4�ɓ��Q��_���v��^����q?*�se�{�9Hr�nNN�������h��(���2�f5bi)����ӡ�:�-���=�:�'t��b�ER����&+)��4�w�<-�����J������4��6(	~�K�z'�0�xV�|��0��ߩy/�W��)����lx�-7�)��W�CNA����[�J^�M��z�7:A���{�� e$���"�	e"�U*�e�`/��Ao@y���R"��p�}�s���U���Z1�z�~����lC�ߘH���<q͞42�a%
���\���K�*ʃ��/��!Q�Y�6��H�����r�btt4��P#��b��Vu�	��>S����B���6b�|��E�n��V����ٶ5"�M��(ߓ���[+������J���� ѐ�ds�=�En���O�R����=N�M�j	���a��L�"��` ���3�l^���q[��В��~�Z* �߉�8�H��_+m"�R�6�@������ݒ("���H�&�-����@8��{=����{��0O�,�ۂ�KFAI�O.��#�}�y���t0�|�	��cz�}��z��Aj������bo�f	�c�}j�����ݹs�SO�gch �c{�E�to�DG$�*��K54j˯��@3�Y�L_�$ю�^�)��NC������%%�<����A<rj�-��p�P|	b�\�ٶ/K#8@��Y,��de��4*Uj�T�#����^�����sYд����͹�NL���3uĩ��<(ȏ��(�U�𮯡ۇ��%���f�T"��T��?[ZZ�ӟ?�B!���0��Y���@e~�����8Y�Zֳ�,355�s�
2�T�
�-�pY:Z�ϐ~��@�f@wg�v~^� h�<�Gg��K�e��T�8��y���S�L�E|!��v�~�2i-7�A�p��\�KLg�޽w�x-�ȟAЬ���i�B��"�J6��*�S����ZE���ǥVQQQ|�h%�R/��l��+55;X�K< ㋷�~���:&0�<��/�n��d�_�)(�-�J%)�1\H�V�l���MO�R`�����h!Y�������|#� �������^��JK�E�%���n�Y��f�A.Nd��!j��m�u?��g��� mHP�H���f�eA���i�[g���Ql��S��G�do9��\@J����뻻�>:1R`��7����R`��^Na$�F�/��X�����N#ᴸ'�LBw+�C*I�6f*��R>:����G��S�H ����������<k�^�nb�:����S�ՊW���Y��ô�u�ʴ��QJS ��KCf���$T	`h4�[?L�:w��T&������#�����
���fdNy���)W^�\�:x�H�'��Ǣ��B/��{�&Q�`���&�gym�5�~�'�z}����5�����p��O�����lT�^��ߓ���̿s��˷Z:�L��4"V�W�Ł~ о����UG�1؄T��S{����N��J�Ԫ�]��'�@酻*�؊q����?�'hO�,F)W��Zn���9=��4K����)��#YvL�0����V��%�C��y�g���ǝ��� �XE��suz!�]Q8�~=V"lh�mo�a>�$�� ��m[�hQޝ-����;��)�cǎ�I�v����p+!(<���P�>��i��n���s�N�V��pJ���.�$�@v)�"U�����!�1��?rf��5L4y��@Q�p�"n~l*\p�[iEx,z ?��<X"�\�;v�rp�f/�y�T��O{�����u��)+=|`�;u��H�9�E����ǈ��̋�6���1Gz������z���as��B1d.SWGgBj+��$+�?����T�������|;�R��[���˃��X����#}���u���W}��6O���5���3�C#r�����(E�Y�5��vpY�&i���OS�+R��w,������6��g�\��4�R��)��Ν;_����X�C�u���ʒǎ�N���S��a����@u0����P#�6�oB,�Qi�o�4 xu-�f�T�Q�hOQ��L��~#�ߞ�i����3,\����]-��&S}\Q�Ͻ܅Z���haG4�~HS����Y����f�eܜu�Im%i1�©���9�RiF #��ã�Ux��&���2�@�^�
�y{@T	�7C����>�#ӆ	���<l�z ����ܢ�9��N�[�'���=��R�8̿�Bf������(��
|�?9[�7J���j�T�3?;F&tnv�	h,�/�[��%��� q��;�;�<\#���QH�'N���36.3���Q����v�NUL+�t�:h�f�\���.S~�"��A�]�[��g6�FG`�#�'m@���}󺛑F^˺�����ss�Zr���U�c��@;]?YV���p�(/�X��� ��'�ɐɃ�*��9��@y�9���iu�Z'm���5< �٠0��a��@&jb���D��X��$��yo������1�s\E�2!
��~v>H1_��Mَ������rN'c�Ϲ���v��b� ����D6<hx�9�ďM�k�T������TL^�����|����ن�C��/{o���B3��
)|:�'������R(M�T�7,!�@�Dy�ܤ6�%�m:��\���,]��Q�;��z�|$�4Z�Sy��?��v刃�ٖa��i)NI�f�Q@��7���
Ӓ��x��)����~Z�j�:0�*��6Ee*�AAQqG�
deY�DA��j�4aɰ��(� K�,���w�r�������3�w��C_ov��1j����F�7���?4�J!E�
�^ǣCW����!�Ą�ҹR�/�k,8��o=G�[J��	��3����)�3}���}fUku��M_�p|\��=�%u,�c]Gkkk9�����AR�/ى��Q�MaRRXVRVfq_��n��Dg���anV:p#��w���e�M��Ōҋ\U�#z�\zh��Ǒ��=����g=���5P�l������	�g({�:�s�T_PA�Z��Bk����dp�����|wq!��Ǧ�#��5�?N�IS�8��0�Xy��{���\��s�[�g5�^⠅��6nV�jv�mX�(�x���\���#�������ǙuO@�WY���t�����e�n�f�� Eދ;>��K�y�C��� ��*'��s���P��E}�VnZ�5ZI��fY�s޻wo�@������}�?`:9ސ��t�޽�cy��I���?�s)��ܺt��/e����x��/\͝hD��9uy�����l��Ӟ�n{[���&SZ�s�����ㅀ��S�}6Z�!L��t`��t�vIFg4� , ��;��!@�:���r=2��xK��)3e#��i��ɂ�.�u|m1;;��4d䩅��+F����^3<6�������傕�5io��G���b�r(`�j	��Q��L�5Y���w���x��}�&¸t�̕���줾��] aT`p.=gc���vP�i�z�ܹ�{��>Ҳ0���Mj�ճ8��;ǜ={<�ѿ�����^h5'�ɚT�GsȀ�I��]�6U�Wj�����R�{wd/��<�@�G��g+�b6��*���o޼�B���V����" �X�y?źf�Kt+�f���>���т���w�)���K��#�u��8ٵ�<3Ea�.c4��[1d�|����U�cGM<�L��������n[mq���K�c�x�N��/h�=�I�P_�F*A����^�;d��f�MH��Iofһ��Z5?��3��_vLA�<�>{}u���%�θ�k�Wo����a�f%$h3�,�-Gx�P^���+D��#�^�w�Y��^*&"����TR�Ϳ$�n�u�3���P����F��K=�0��l���2:ԛ�M1�Ը��P���y ���0���֞�~<ߟǷ \�x�9C#������v�in%�?��ry<[�Zv�H�:2��?"���>Wa���qH������_��.![��٘0mu9}��]9��l^� � T�;a`�t+�t�l�B�s$��ߨq%�粓�<VR�vU���q6ױj�������[{��1שJ	�"H���1f�2�-�dXE�{C���	��򢷇��S�qZ0�ʺn��		
���:*� J�i]:`&�l���e�{W�1����?�]-\����Nj�Ff�C �*�`y0N�D�����nb]}L���hŀs�@*��:���߄�5}n%�v^��f�#j���B��}ł��ʲ]��1u����u/�&" �Kr"��Oѱ����<�=�fy��F��\�)����e��z���]Kv,�#��d_��`��
��,`�&J��8�߭�g�?��ӈ����B��^S}޿�j�,��$M�ka�S{���m�u�=�@�M�Z��4����)N[�\���F�%��}� �:��l���@�t�: ʤ��a�H��0��_��,܋aC6,X�[-�+��p�O�l�6�.<@�#me�IHxϭ�O���h��9@���ѐ��2Cn�Y����b�!gT;�P}��dY꽒�����.�~%�%i� u��TQ�~l[6�Y� ���GaŒ�{�����
�Gv�Q��mY�<���T�{)e�A����n���MK���nX\	��w���f�MZ��޽�4j���utܵ��/;��MG��Ka���>W�o��B?�ҭV_�.9����?M-޼��}�Ϝ��W[_�:k��)k���s+����By�[��۶�¬�?���l��fz� o���7|�����|Y��*nȻwʮ�׫�v��<~�5W�ox�CB�Z\i[[��D����|�f(��j�P�6��*Ca�&�*ԫ����ȍLG�l��4���[�y��־�	���/Ճ�c��|>�~d�s���J��X^dN�b��s���0!��P�HYc޼y��!j�� ����Q_f��QZ��]qs���ن�����f���Xu�ج�*⪪����^���d^s�ݳ�ɥ����2��6yp�nvke����'�����U�r�8�gb+�a���D]m����13739��:�8K��ϒ^7��.��9 ���5���#;�!���t���?����,omjXɴ����I���@-2�X�qʝ�� ś��k}����
�Z�^�\r��ms�^^jjW
�U'����Q�Za���ɸYI���U��s�����hů�~H�;H�������ޡ�pt4&�}C����+AS72�}.��B�ǭ�R
����c �^;PYӌ7U������DJ��F��G�k2�����ϐr�[f��t�1$�y&��>��S@�be�����ݟ�*S��:�fGj{5��Ǐc�mթ���&O�AH~(//_���#{�)璲�'��IN�[˘a����S��0���!��G�����|������] zl(+�ml���@sP�?�ĭV�?��ƄS���=��Fx���g���D_T����)L��r7��X��<i�-X��X���X� ��j���:��Xpa]�C��t#�����i�'���~yx�#\:�|}G��6��5�k�ɓ'W(#N'�n#B\�M����2m�z�ii�1E�el��~@"�0��������ξc��vWG(��Y���ř��7�%sY�Q��UX�?g�(��6�Uc���{ۈ��&�v,�u�%�����b"��&_/{482������3b��f&
F��\����w�%����P�����6>��%+�z~�,�$١Ƙ3g�z�	SXk�v��z�wO���8�"�Zq�~3�ʹ 2J��'��r�X�%w;-��P�6e+5����>���Tzk~�޽�0Ʋ�@iA���K�g҇����bw��\p��?�j��Q�d���+L�s|lǳ�m��}��R-s�[񈾩Dx���c}(���Gg='M���'�̭?e��(}��<�=ɷ�τ�z�|���=�Q�^gѓ��ȢR<�|r����~�X�Xga���6�N���U�X����V̍�b'cQ��]�w��1l���A>
W��+���1Vw)#�"&(��j���Ȍ<V1ŝ}��s7��S�l��u�SQQi��!�!W�^rH'��r�lʄ����l#TfLv�G[�Z����B�	ǽ��s~�����4�Y��d������&�j�n6	!�?�q�ܹ!1��8X�^�>q��! �2�kb��D<��0n`��V�6'�����O"4�w�q5�p��o�7V-���d��q^>��_��W����ɹ�/8���e)[g�k��q��]�x�bU%e����nL<چh����Y�s��m��|��3���s��5���`e_�� R]�(ɰ���5�����x�s��u�L|9j�m��k�ǭ��5"��^�Z��ו�V��E�h�/��>E5w��}/�5��. �B�j6�Eg��\���/WwՈ�))��Ʌ���?�Q>�E)+[��
cR��?>�zZ��n˱ts��0��F�r�X,�RS�YN�Jl-��G�=k���1���K�c?'W�:��yO��%�c���V|ށZ �1f�/N��x��8���L�q��3_(>y�孅&��3�u��SBe7�h�{�%y�������"tkx2N{d~(��sR��=G��ID�v�4�r�����lǗ昃\���Bz~L�:˖_���T���*'�[���$�C�����eDEJc郗�b�}��$���#�W<���k�XB� ����`�K����^�.����Q:���M�[�&�T�,�����~���U[o������Yqqq:'y����ku�	�2���=#�)z��l"!�"*�O`\oqnΪ�:�۸��Y�����@O�����+11��1�	4���B+ԧ�S��֬×Ń�f,��`#wvivY@(�F�c��z�/�xs:h&Ke�ps���$���e����>F���B)0Dq��atC����F�"K]YK\)I�j�Id�MW�l���7�*������_X�nxx�!"/��=��K���f��[��6l
�6�q���Jɷ8ڤ����o�Va�G�r+�r}��=�M���,�i����
��Ul����A ��l��Pl�g+4���9_ӁX�B�$v}�ZG9��Y5�hk���2��N�L�n~�=`�F����\J����e4�S3��9����D����8��4
R��֥\�������q�T@ů(&[�̖Bo��^�P�ۀA�O69�V�v6�]c�*1�"p��ڐQk�����%��hA<�}���E����L�h��@��0,꾥����+&��� ���u&L��$K�b�B'�%'"X
�oː��`<�!�T���W��u�A+�	B��<b]�d��VF�Az�e���-Jr���jʼ爪s�	��o�?oE���9�)?A��_�4v� �w�jߤH���c�X�q�\"�?�
:=$X�u�]���1���1�%�r��.{�H�-��w:�P�b�-�ލ7���/.���ת�M9�U��=gR�
1�cm�sZ��"?%T����D����rO,�(��,�z�h7����"	�MA%�����M�=����oH���t'MpZ�z��w=NH&��N�ژq���O�ѳ��ϯ��ɩ�O?��ƛ2x���^&#7QI�B_�4Xss��A/�@c�'M���c��5(��E4�*_����/����jb�:�7o���*6��5uZ�9߂�cʚ�X�y2�ܥd�GYǄ��i"�5c,�9zכ�_!_���[�Զ���?A��d����F��x�gr=��?�Q4)��.�V	����ty�)Z=e6��*=����V`�1��� ��)P�@�z�-��.ct=.��2�ɓ"Ui�7�ڤch�[
NOҘ���%���d�t����u��h�� -���b�#�wd��U��M�x��XA�ܓ�]��75�ɜ5셾�*��>��Fx��|B�ƂӪU�@n�k����h�Ն嘠:$AY,h����W�M(��C3���-	�ύ��'%'[̒������$>��*���x��@��퇥�qm�:�p�2�hy%R�[@�:��F�[c�J*P�ʔ�e��3������(!.dܘMO��f��h\�`9��4���	ǧ�������|�;D4D�.�st�����M���I�r�ZO��H��m�33�m��H1�ܸ��^�x0�[����J ��X5T����_�K�gүnuQku_�5����>W/�4b[���F�3�̝|��vE@]�qՍ7�7�=0)���e����c�*�t��<���^:jz����y�k��bo��W>����/w(79�S�C`ͤ�������56����������=!K�x���Z�w�o�L�~����P��hR<�i��Q��F|+,�믿b6�N rU��f�4E�c@D���P�R�]��L�	u�q��j�ف���ٳ�]8�d%�b��4;�wS���Q)ӡͯohwW��c�^��f�=��感sQ!�I���������������R6�������_Ϡ}�_�M_�1�Xԏ�o�ba{ �	z��(� �$)A��7[vlCK�7�����G�TVV~ĺn|�h?c��Z�sv�ЗN$�)*Z@+�.���*ӏ)8���;�<�y� 	o���@�6�O��>�%%3����&���ك�c����$�������U��
�FXJ#��r$����|�
_u�Q�Q1;9'+�ݝF��o�P���(�����2�|�U�'05��遁�J��P��照\\>��0�˳���U3���d(Gs�y�P�g� %Hq���$��Zn�\��!�!���v��Vj�`x�͟�4�n���d73V������i��j7`�h���.iZR� ��
���H�mA)B��u�g�r�= ���C5�i���,E˗->��k����Ѱ��'�bhG1�*٪��dܙ=�9�7m��E�?Kz�����N����cyFaaa���$���z%���  R�J�\���`1.A,E����飉�5d^��@�wQA�[����8=��ö�9�u9}Kq����p���f4� ϗ�� �|����y�UW�#Vg�&����;ȗH��5M���Eˇ�7�&?ߥ���%�8��PJO]�~���W�\H�-�2u���78��N4���fՊ����ki|��8GU׻�Q�0&R̎��X�0G1��C���.� ��JVp������9���pw|��9$y�7�-����|�X��`E=�8�"��>9��j0�,�Ӛ%��@>���A�Y��-%++�&��I��fn�,�A�A��rٓ�%�J2	��a5uS���Ji��h�Ϳ�d�� "��`]�xJ��2-7�ŉjkk�}�ҋޅu��N�ڙ��P����qf �#�����=������
]�N>ٶ䪡 ��W�&l�ީ��f�ٔ\�t���
;Ŗ��$��ݑ��}�gZ �i�D跋�s�U��s�Фxu��O��������\Z����{nC?]�ZO���Qs�i9�Gc7�'���$�L�#�����e�޲�S�g�}ǣr�@�rr�
zY�%�Z3��8dk�C��[��E>,WU��wb�~�N&�#^��o�u횗>kx+Z����޾�> b�kB)uL}�<��Ј���I�N�/�		�6��^x�;�#u��CG�{���3�-!�:�P�Q��|���P�������[(�*"�c$^G�1��q� ����Pw������?RRtv������Pr6F�\ �D�� �w�c��%=l�u��U�q|�YӰ*�^=J�>�%�h��}�@��)Q<x��C�����_s�2 ���s�|=MxLn4�s=}p���ӈ:�=rlI3�ʌn���Ŏ��M����I:Zo�|X����0+�ˉuOr�S�M�����z���t�!��.��.�����b?"�-�I��i��q��	�qTS�]���F,cw:�T�2��Q/tV�vq@#���V�
�5B���j-�7�ɚ���}C~3�����?O� |)���7Ѐ��{����y� �����/3`�{)~�A�儘2�y,O���r�${E��[W0h�U߁����x}v����g�(�n��&��\�`���jw��i@x݄�"�Z��cT��J��j.'�k�
�������Ƚ� '�}���<R��{�U?�u�@T��K�����(L�\�]�+�٬ex%��؈�Ox�4���s���,/���KӫG$��7�m<��Xڰ���8�P�����D�KG �۪S��D�ϡDI��%�y)ѹ����⌀���zW!��٭���z�XT	��!s�y�M��0�����\`���^U�A��5�-#~���0� ����y���K�q�oA��?��j� `���Q�J�@�A��1<7d
*Zt�2F�����c�d���ʠ�n
lNms��6'�UԚ:uj��;��d�{���G����_�q�e\�a0���-?d!��cµ�z���C�|=ߨ�k�o
bL�^��T��kwo8���rQ���_��0)��-���b[�BM.E=T�g��W2��!N�]�y�&�PF�'���	�yO�YQ����\�L��|����nj��f١�K�x��u�Q����ܔ P�����΄�� b��l��x8ڦ(L�tj��^j�����pQ�����=��#@���Y˅�n�d�vv�?0�G�J�y/=)1�b�2c~�m��k>�;bbߝi&E��?���Bk�(X������#���]�Q��u���߬G����sKp�{�ă�8D\��S�)����>V��f}�k+��-s��#PC?���c�#1�X�T^� Рq�r�<Iϗw�5���`��=�s���_�D�pM@�}�;�;����B�U��{�%��% \ރMixنl��"����֯c��B�7_���
-(�������C�$������X%b�!Sa���E��>�a?�I�"��th�jh�Z)>g����紧,Ƕ��(0��|I�ҙ�z��uV�7~s����nfZ]����3Sܸ�����=Z����1������;�K�҇����k#}răg�������]�0v�%�zI����X��&��X�&>��h��p=�t�0I|r��6yT�j� 9�R`�Đ�g�A�=��[O���gCX�9�ܖ��<0����r�z�:h�����X�x��%!���I�KC�Н��O����,�q{|�~�&;�i��g�+��\o���2|��j[�Pd*��$�$��80���?�
�ί�H�'���W2�Q��Z���>(��s&�p8�6C�&d�A[�45��CeZF�4�^���\���e��a!H!�4l�z"=-�A��$#��?�j�,S�`�|ve³��B�i-�����A,��3�M��o�mV� ���J��V�Q"�q��zL��������/I�������
]E:��[F/���!2a�ؑ�G_	����CPR��1��'�2 �7��H)D	�&����G_$��`�;�wX��? �6fP��L8���*����������G�����Hv�Ü$� �ig�62��{@��,��@�}����<�������[u-�R��Lg�����6�|��w٭-]�$���Jzc�,Z�7�'Bܛ0�Roo�� �\�`���8F/�6��MUn#GR=1�K |�8jc�����P8:�� 5��;�+�g��yCW�~.��18��XҚ�p����苮@�8�F(q�Y��BSz
��qC_����766����]V�����a&�Ka����"W@�qiii���}�OU�%W���聀���"# *hqޣ���kt'����a=�<�Q��u���~{|>w�Y�L�!��E=&œ�Nx��x����:^b�(�͕
�\���AZF��b�y1�i���cJR�qKvR��j���Zu�eh7R%h?����9/F�7V�+�8L��H+X,���J�u;��x�DQ�h�y̬��˝�ܴ@��;6L,� )_�״U	��4E�y}����gF�@����6	"��h˶R6W
��Φ=����eR���(kV}Ύ���zտ��hjz.c�^�M:��5�G��Ϡ��@͂"��_����6(NЧ�|[�~>=����,���J�~?�z�N~�	���)�͊���>º��ݤß�r�4J+��U�LE���Ķn��i�x@a��E�U��ڿ�rl����a̐e�F��iP*s���Z��ߨ-_�Y�č?]n�ә�I9��s- 7��ʊ+�_���K��9S�[(�?�I����5p��S�Xd�Y󯉵�_Y�ڀo�5�&qBޥ[Z�]�vt�a�ŭ��~Ox����b��åf0/�ا���p6��[�a|�� �Ԏ�XS�	�f-+!���dO���R$�m�[��:��XުG���*�J,�W=�!���A{g���]�-�K:6�F���Q�?���������c8�����Ol|�3�����!��3Q[��bd��
�Kp���Ƭ��Y��PK    {�X�?HU!  B#  /   images/585092fd-6de4-462f-8499-92296fb2c536.png�U�S��]:��n���	i�F�;�F:�����n���n�x����	�;s�ܹ����=s�<��@lJl   TT���� $lL��m�����EA� ���o#��hB�]R���u�~�t�0q� xxx��8ڹ��|����l�y*A	 0�+ʂ5=�N�<5g��=k�K��"3c�����s�zhj>����v8�*����U�]635����D2a���Dc������M�P~��"z3����l�Μ�ws�+<����1v��2nh���0�*�� �dz�̗.�`;7)�G�fK{�"j�R��6G��e��o���<��Z��o5І�h��+u�8oi~�'�f;- C9p�]t���F�,��0^M1��D�K��7T��*��F&���Jb��{.����a���"�P�R�9)��H��G��3qx�N��
����=��Sp�IP���=YQ#��Q-��\F�A� /R}cЩs�@} 1���H%��4�k��(6K
w�Uxt��c��[?2
��Gh 6P_�-���(�QXA1��+6o����ws��p�&E�{�Y�X��"�UPӊr�K��=1��8��K�K o��H�hV����[9�p~S��}wuZC�p=3��GPZ�d��-��jn7��~�ʸ���O�֜�����3iZ]2nT�p�'/��g�}�iU*�k�u��V��gOaG���:p�r�N�@��^\��	^������N��ś���4��Q���S��g�S4O_��&�\k����ീ�A촱4��N��u3k&lE�&K��q!� C؁HsCY��ۆ�@�[<�I����|�h5�@w��6�:<��#�w�\�ն�iI�m��G������,�}�f�ԁq�cc}�zu���'�4�6@[�KW���<��T����4.IōˍY�*��1�ف�+���R	^��>�]Ư�;W��d���tV5��C�xłyx�^hE�윽���d���7��7�S�+tP2�]��1��E�9��j����60��Aʗ}�e��3�vi#�k�cNv���� M�U����D�@E���y�̴o�U�;�]�t��n(-�"�B�}�2v?e���}�;�{��'��{�A�/7J�3�f�#��{2���t7�0����-��'@~z������
 K[���ϗYSIܯ�K�>���@ �p�^��z�k�w}�}���f�,��sT�yzU͑6�3s�7G@k��1u���ˀ�k7��q�������������>տ^���� ݔƥC��,U:V��3]�u�������&C��j!���W�>ȹ���/be\~Ii
�l+�����`$E����Χ�"����O*������|䢤W����'mo����
��glFE��_$�)�xK�EC�~H"/לiVcƁ.��4��tFNX�/��Z�3���Tlڶ��đ�Q�"F�VV��ե<_Z��������X�>��ADr�_��-��2�M��[���Y�£����R�"����R����}�$�b�E��x�@#���H>g� B�ӆ�z��F�\��@tR�>��d���9�����8������N�1~��Յ�ly�H*�n(�d5��cؑLG�s3����j=m��� 0��R�ˋT�eM�-֨�B.u&o]��?,��aGYA��i�L�s�x!�5�7�������hpy*-�l�_�FӹaQB��s��c��ٍ��4?��\�uO��`�j�!�����|*����P�嵙�1�@m�º�t�:���g(�<g�3�=��u&?�[GG �ڗ���#�ڐ4�Я)ٯ.���wޅ����0����(-�A����yC�>[}5||���[�
}	~�6T�J���9��x�x�4DE�|��_.�1�.��l�6�Gtj��;o}B��@�����̛��/R��J�q
!3�j0���[@2���}8Cv��\�MV�iM�(�L���� �G/�~S�߳����������~"���
������ߋ5�yW�O�c�2|*��[���3j.-��ބ�"���rmʅ��m����߈dd��$NQP���f�546	{���|wRZ�I)/��Pάk$�3�6����~�RfU������u�ס��R��tT�6�u��S#����zd��y�w^�Y��E�'�����H`��i�1�"+�ˍW����	��W��0r䳒s~�tC��5�n�kZ:f-��j�7��g�q����7��#M|�<����
�梕ѭ����+�E}#
�̸sૃQ�z�� Q[o�伿��:!�ޗ�qꏳL���XY��p;~��~���ΩEMBD�sw�M�!-�j8�Y��dT��k���4	����c�*[��P�4�4�.����
�o���� ����x��t��������ye�o+w��T�g��}c�;�#<�H�<geζ�����_S��R��5pVSP��{���p��7�n��P��<)�ͷH:��uj�RAҦ�(�����ݳ��/eB=�g=v�	�U���62#]75Gd��nt|l��s+��hfn�ɥ�M�N�Om�"�aTF�'?֖旱.��|H"�ǚ����ϛ�>lس�r��L���޷7	!�`US=�>4�煖W�FNú��(q�asǟ�Tc��6P����Ie���1�S"��T.���n7u!�f4����os{kW����/w*�����.��%&�b>�p%�ݾ�%ߌ���W�'����q���O�Qf�B��!n8�sn
�~j~���|7�VU�Wj;CH��99��v��\QA���o�;�S�lj�٪V��Wf4��H2�8��د38�T����ėh#�f[����M@�E�'4�Yu޹�������e��7�e�ٞ�2v�+���?=��9)��Q�#�S=Bxo�k�0֔��2��l�M'}��B�r_�f��{�7~�W����<|KD��-C�4��Uʼ�jHa�
m����ث8��N\����ZS���Vڋ��G���瞾��l��zn����'��l;�W�m�K8G	���[��?�c>H���J0�c�����;�?��w�6g��2��(�1AQ���M�y���[�d��T@�i�-����X[X�B���f�0G�k�d�_��7w���1F<�l]�>�^��M�	��q����H�KzmY�82�#�s廛��E>.&�۳�ǥ�g0c&,h���6u*����U!��2J�|^Q����9:gr�x����]-�*o�F�̱�`��E�@�Jho1N�2[�^S���Zf�:?�t���T�Řl!\X�����
�0hP�"�w{ɭ��RiDc ;a8Ir���f�[��}�o"P�'��OG&$~��4��|nj�2��oǺ��Ye��!�<?��KY�:5�+f
���ɡ�8��\����L�����/
G�C��Բ�9%vJ������X������E���7VR/A*��sBN`L�p9#�(�9���c�J 9�O����FOY��a��k�IƘ�����BpBSLI�*׷�G&��gL�a��J� .�rǥ�6�.v�_mO{拃��~_�,�a��y6��@��4m�\6���B_�	L�𣖏���g�֜疸�TüO}�>�㇁���������>��	o<ƍ�������>�x3���H��Z;�)x��t���v��h䏲�Ws��ѣM�JgBSW׻/{=�6Y�/}�G�a�|Tၸ[3��9ހD�)l��?M�7�\ա��6���]fq�;�|�0@	�/L�IZS^|�a%��Vz�����9i���G���﷞�;5o��.p����7�X`GD`t>�-�Y���0��o���h�p3��r��;z�q�����B���^�����`�vH�%�%ͭv(x��X}�c;����}`����H��yL>0�`��m���[0g��W�� )Fr�Sf�$m[Kx��z�	�۫�G%�R�O��
J��+��F�]v4�9���;I����L���8��ҍ���wN)i1j���c�T&�M"l�"��L7�7���)=\� ����z�g�a��L*t�jB�g'�:2���������2Оt�raȧR��y����8��YP�Oh���a$6�!8n����,?��C'���.�M��#����nj� �~��K�nA�;�k�u�/@G�]S(�<k�lZ��Go��Ϊ��\c�e%�d��k�1i�"�5� ��=��t?���@��ƕ�8v���wE�Y������h*����r:Ɯ?�ms����l�Rx���~���o����~�F	�cں�?�Q�U
!t�����mEE�5qs��u���2�Y���-IJ���<��&�KC�B2���ʀ�]~*IQ�%.�Q>9w+3�@^�L]���`@X4���r�Æ{2�`)��<>nLʾ�Bk0<;���yK����ޘ�J5�A����n������HƗkh�K	�%,�û��Y�K�>�b����T�֓�P� � �ΨR�V���fM�{��;/q,T ���5m��'3��6s�׼o���a�֯b-x�#��}�q�Kv�7i�O��R?@Ӣp���/'e޺"�X��ɏ�����	-�*�p%����A���
�����?��nD��@�\�f�t���7n������XϘ��h_I�ˣ�1!^hf|�VS����.�'+�?߀>��^AP�fg��w��1!蘧qs�����xAp?�Ы�㽋��`z����6�'���f:�8��l@�
˺R��l�@<*���h7�Z���<Xy�{�#���L%�v'S~W��z��T9O���gc���k�U3�@�#���U�z����WAV����S��om�:Gx����U���xEf��b�J��:��,�D���������_��a��N�(����ο^^2l����j]�������#��Z,��^t�x��&x����%�A�9W�"�{~v}����t.�����H��$�h[o_#�fá�<�,��X?hr�x�IȮPJ�n�w�����d�&�(x��L�����K��^�BQ��lc-$����mog��v��>F���}�|�S}g(n�y,�\e��C}uv�i.u�����~Rm�*��MÀ[�9Va�/��T�ę�M��0�fz�ȁ�����E<��??��3�N�+fk%�5z
?�#f�(�*�����z��'�EH�
�:pơ���3tL-�?� ףg�Y	�h�wq3�wY��Ë�R\�d�{�����c{|���㄂<����/S��Y���f������,��C_�Y���Sm���ay��.cy`�n�͘����!Z*L݌����63�us3ˣ�c ��ݵ�h�~C%�A-�.�&��`Ƀi�U�H�*�~r,��i�'a����ӂ�����k,eFJ�`w�5o+���D|d�ɰ�KP��d�:M�`q��~���H�@K�y��@� �cidf�_�=c��`�b�yJ��-O�8k}��b}x@���Qr�bIi�\P3��,�a�!�_s�����K<����v�y;��j�WU�4 {��}N�b��&�$dL8�[c
������*�ܙ�8�B#F4�F$��*�~ᚾ>�IL��D\��7�6y�lHY�E��C)3%�᝶�nzl��ë&�G�$&Փ�B���'�`l *#��͙G��i�7dij�ߟ36�Fs��e
��xW�<Jj�i�y��꣰`\�H��b$����;�c�V��DRŷ	��\U��ͭ��y�آÚ,x�{��K��R?��E %�GU���:i�@Z�H�������٥�o�r������p��9m84!��9��q�P;���c������q�N���`�<�_m�_-�O�}�w\�N�Z6���ƾ�M��՞�������Dٙ�b/�BW�M�XT�8�y�����8CKі���8�h���T/\T
O�Z�V�L=��x���,��x�v����J%D�����i��[]^,��G�����>z�I1�E����'[�4kq����((fܒk�x�`�9�Ń�7⏑�Z/t1�$W���{�t��s���ܠ�UO�s"i���'�X3���>2�������O��j�#�]!���IhJ�D<]���������I�81��2��6�|q�iǂ<���Nr��;9w�=������8,�X�&p`	��9w\
VG.�8.q�EM�iY���@��q�1m�j߅6�}�	��Q��su��`�w�Q�i�[�l�!fg�>��m���wM$D^��+|>:��˖ޫ��Yߝ.6K�=0č�ө��e���h�s�{���x\��Y���*�f����\r.�
DQy:���[t(5�jM���d$���K� l#5�wǐ!��ɿ��Y��D*��;!��!9�wŲ)��
]�Q	�ֿ�/��q���������!H6���U�o>1��A*CP|�g����)v�J�������~A.-�rE�6.�(����$.���H�)�#t�U��+� �G����_��?���/�~��fO��)|rn~���S�Fo�7���R5��|���:�?N�d��b���g*-J�[�'ʺΝ�V���0��KӠ��K&H�'�������V����!��rC����ڳ˸��|5i�r$KȳA$��r�h�P�-T�'z�g��@�H`�;�<)�E�>��%^�H�6����n�����M���r�\�h}�*��V�4��Q�	����G������AR�M��G!N����v/0�����zy�����Q�!�WNqY
��o�04m�[�9�qQp��o�W�fSB(Ku��#�<'��'ϭ��gB�_0pA�bٝݪW�FX�l��I��N���2�&�?�����0(�P����=]D[�>302lv��̫��<⍌�^¤��q�Z�О���Jі�H�⿷~��[>�U�R lļ�R$y��!*�(ǻa@}Ne��`&<�!�I�ʐ���ć��m����+�&@�E'Hz9b�o&�R���&-�v�hyA��<�}B���Ҥg�(�!�%�jCP!G�jNnnD���ژd���.Π�i�U7L����\[���	.����!�A�{ Q�Y��?m��ak��f�1.00�S��!�sSA��f�%�Np��(�����-<��t�d ��0���	j�$L;j��
�\�p���ڱ�������{#8�x�ˌjN�TnU��f4��u�o�9�uD����F<R��e~�>�Kb���$3���D��x�漹��h��x4��a@������_Fc-�(��7���O h?��~I+6�~��/���h�Y�i��_�A	�������eT�$Ўl�U�3:
U:�P��W�6=��8K�V��7yѰ�*��$C�O�d�J�D-��M�S>EKN�*%Y9*�B絥���*7'n�JI`�CFʄ�w�����	C�:�.WP��1%�3	�[�lC�V��G�;�h�Pd��]4G���P��l4�=@��2����?�#N��µ��F��!_�Sm�4����dY���+w��V�r;�Ovd=X�~ɠd�3(,�WtL�jG|��/�B>�Gi}%聖3�1�T`~�#$���I��a��AN�'���,|bHM�3�-�"_�_4��1|���P��8E����,�@J��X*[)<߁�2���r��B�¼#�a�=�%ە��A�Wߝݷ8�^F7�fz��R�b�M�n-�k�A��\t��_P՜~f�MG'�sg������Rn�7�Ѻ����"��6�5�;(���~A�nԹ�
���s��6ݑ�����Z&� ���c�I�y�?�l����ђA$�͟��9ȧ���f��cPUg��	(u�>#
㏾��	gA̡ɁX΄ZcX.砮���hT~Q�v�z#���ph��'7��Z��Y��Z"��Y���b��p��2�s����hS5/W���G�h
=�=ZY5'���4��3�����WY'�����,Cf����d�:���*���#�W%��W�x�s��_U�I�홗�����1\)�e�Er,s5�r��YH�H�q�1û��@2D�R6���
�6y`jWDA2+9���Kf�L��9l.LU��v.�@�����x����X��񪼗c��`2�(	�N/΁����΃B�,��F9S8m[����Jq[�07w,+��
zE>�M@}����V� K�ZspK�	�щ����M݈�D�-MiuQ�|g�9{ٝ��|�C�o�k�n��Xdy*@��*m�����R�g�1R-Ks���9�d��j=s1�m��x�sms�O�1��[��Te+!�A�PK    {�Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK    {�X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK    {�X��Xc_@ �d /   images/a9ae5602-6322-48a1-b803-2efd75c9b3bb.pngL�TT��=|))		)iZ�D��P�1()i��a�:D�{��B��;|����]��r8��'����c�kUyB|*|  d4  g ������ۤ=����RQ����E��N
�� @ۊ��j���?�t��s�t�rq7�`	���s�:@��͜,�?X��R =�(#�呺5��=���z�&n}���͸��{�����V�����lm'�alɾ�#~�������r�8�X������sk*�yg`���l����E��{cg^�ă�z��ݓ���� P/�޳><�D�I�)�n�jw͋���5�?'1b	�R�+��9Ϡ�l������s^_�K�M�{�%U(m������
;?Ԁ���?��2L#�D��1���d��	��rCv�#��}�)����(N\���x��O���_DҞ�`$�p4�l��������M�}WJ��&n��G��8��3�(t���5*z,  ��$F��ha�.B=F�'���\�Ϫ����#w���o�C,"~o5��Q+����L��-f�#�\��⥅V�t� ��H��A����W\0k.)7X�:(z[lq�� �.��M�z.'<�=jC���:�S4a����7�M)kNk�y� $ ��8J�̵�rĚ��`��f�Z�S��	pw��q�J���\�m���T֥�\���읮`T"�\vE��r����ӳ����y5;�ٞ��� ������V��[LKi�G�L��8 ����n�L؅��%��
=��np8i� ,�ျU��n{dl�B�����0o�y�*���=�o��������n)��R�:����O��;B%Uen��U���u(�3GD��@A����9R���uy@n��^�r��B1�Cul���b,�R��侇TazɩTU�:����ĢQ[���3� ���p�x:�����������m�؅��N)�����J=��pd�&��U� �Hn���6����4+_~Y��yu�`z��T��&[Ѧy��ü�Er� E|�g�9{�&y��m;��bTc��!�u�(��9ucZ>���;@�����p�j�A�6�یt���oRx��N�4N=9�p���y��d���$��̗��#������%sr��,�I+J��E�/�9  �ް���`����k�Q�6�Z��&z�ji���T�U��(lQyp��C�	�եZ̑�m�-DQG^	>�2���O�X�����dY��k�<C�y��J�^�?[�Ґ�8�V"pq��G�����oj6][c[x����3�-��"�r?�c1[?.��XןRceۯ�M�ls%�0i(�/Ќr��n��q��U������]�PHl�H%�3 Ѕ��ʔ����LU����M�T�`ꔯ=�S�m�QI�G"��ـ	�/�R��o5�&B/��'�}�N�ܺG�ֈͯ�() �}�#{��z�E[�t�h���0�����14|��`����jf���A��M}t��HL�v�P��_�Pq�4k�7v�^2��7��kOPפ~�<\5z�N��o �^�,��gvn�6W"�]���kOG�d��y�2��O��oDw8^g�g����ς� �9�͝I +s�u�dh�ږ��#��@S !䠥�
�L\q��-�u+��ݤv�hs��0+�z��dL<�E&ԜӰ1����v�����P/ (E-�Oym-q��o���SZ��Oo��(Uz�YF@��'^R��a�(�s9,_a��&4���b��W�$6�p��C� �d��������������o�&�"�@�TE��anǮ_?S�D�l0-?�c$.�l���k"'m��Y+W��G|���Zv� ����*��$_+���c����L��*>�8Sax��\�
p
l�����\��`�9���l����M]瑳���\֥C�;k�Ɗ)�Rߒ!C����w�c��!�����{d��a�u�X�?�H��H̍�<��=`��KЎ���xH�K�ؚ�H9�����f?���L�0����g �jv�3xb;�j%&%���Q���vp뭔&aݴYˎu�E���G9��M!�s���M0,?���ѻ�yXT��UT$*v;��Ya�m9��]���B���0�N�����W{��0���>p\jpN��&������[x��:��O'�@��Wz��c*my���s��آ3Q-�?qh�K����5�f�Rq���j�g�#Fο�Ǫ����\`�����Z���W�o�o�O�%�;j����b��Q��
�k����+�_E��~L� �n��h��q#v�#0R�B��_oeD�3E���m�T�2��	;��+������໘X�)m��4@2bQ~r����h��۸Px�xؘ�����54玎[��J]�����3gJ�뽀v�,%ظ�w��!�Y����P�� b���z����}l��G���tǲr�����ˈksn�b`����=p��������3Hci�ì���{q�5�r�p�ܓDqpe�����2���i����$j-q4��"x�q��M��'�q�t��X�k�x �DN��P�0;E?�y���@�X�w��xK>\V�ea~i�t���3� 7/@cS���CAc��~��׵���ݺ�]���.$��̍�}5W��|,`֍��IaL�p盽��t��7��9�� ������o���k'���X���$�Ǆr�D[��7�up���H��+9�\?�uLP��῕�O�]2]º���:�U0��SӁIv�u
(%����C[��ٍ�@�l�UA�hI��68���Q�0kQ�(R�D��� V���g��6�D`"�1�~(f���6��{��
�ڔ����t�Ԁۅ:t�P�{5����?�!C���L4�b�a�ӫcz�������s����Lg�F[�_>��zB��fUt�� oհ�[	����ߡp��h��q��|_
��|cŌw�@S^9�.�(޴p7s��@3��Z��4ؙ`ܗR?c��g�&
����U]T����ے'o��+���J�:��7;�zԧA	�inez�y]*��y���=�%-W�?D ��^ʭ:�U�J`�]`��҄p m�&<;��?�n��h[Z�|��ǚ9�B��#���%2�w���ꍛ �D����(�po�����{89Ѵ�eY��� �jq��r67�
9��(g�ad~U�5��� ��n��dJz70o���X�/,�����1(�1{ZS+�eQ`DI�W�^iv�ʝ�s����0�P?t�FsY���4���δ]��G�D��a���C#F4��v\4�ևAV1�t�eJ6��qF��e�]	?�э�<�}����0ۜ�`�ƅ�a��-q	�1;R�e�O<pʾ��G{�2�������H�=?���;P��(Ts��_��-�f�b��&Ĩ8A���;�+-�όK�5ȿ����"!g��!�"���qC��y-�n�����닃�U����*�
��4��z�@�9�ciR�ͭ�K0|�c���uTN��W)�cz:D׶��]a$s��j\D��@4&[����WY{n�!�2S	���S����x;*����s"m��%�3�ꦍ��=�(-Q8�{
�$9�ߴ�5�5?��Y�)X�J\r��v���0�~k\��XO�"ܠ�����4,����K�k��L <�A5�C���6����>�m�q$�~R{$�~�t��F/�%����댔�'�!���= ˟NĞ�ag��Xt�$�g�"�����,��p3_b_q?���];�"��h��#����M����5���2�>A�|im��k��\��x�R����F]�/������
r�!vn~�%<k��)��.�?�u�%��OLe��M�(Q�v�^��p���"Q�7�� �����1'(7�?UP�f��1f��t�9�+\�E���mf����"R~����w�%��UV�9T��Q�_�"��SϼV{�P����D�%�KhEsLO�wO Y"z�ڣ����q���GY����T?�K�*��<j�B�֏�>�
{Dss!3������y~�l�3�A��0-����jXQ~�v]T�6�$�����E���z�tI���U:nT@���5��H�-�X?id���
�5�bP��ՃH�)�#�Ë�/hkW�I)c[:xQG�rL�E@M��;a�ܤ� �e��h�̔�4d��m��g;n�:F�Lt�|T������dAdj4�{������:%�����f��Ĳ�7���x��α��">��F�b6y���5d�ڥ�;X,�fςqׯ�� �����|��J�X6ұ
�<5QR\�lOqDX~Np-\�B  �?�� ��|ԥ��C�1�F��^�G��40����%��L%L�z>�/�_#�i�QU"?1�&�4�s�iQ��Ơ�I}�٤�5�9����"���|���n�3���GRh���:�o˥��˘�epP�-P�,�/�L~��vS���Ȩ�ZDx}��H���L`�2F��A�t�C�k�OE�;�P�������s�w�����:��y��S�f��|l��Q�@x�U���wm{�9�6�|̡4���x
aC�t���=�C�T����%��;t�?��yD�ec/��ۛ�zD��'q�֮)^\�ӆMwn��D�I�\�mm�Nss�"���ux��91�f
�|ÄR-ɯ�U��BV�%d�e��FSA^:�xR�N�i�h��f�0^�"�-�IQ��<.�P�lz�f��t������E.���RK��,?r7�M@�df�k��X�B&��:���N���l�
�}����T/��%U���a,Ԟ�������\� E��T6�4;�{�V��Y�a&��sS9BnB~<?s/���^��o{r'�Y/�����z\ �&�.�Ն�b�e���s�D'{��ޮ��N��z	Hj�5��TB��kላ�����\����_X��
�+.�Zn|�[�W�-P���jH��y��Wm��C�F�^�%�Q��	 Y�\ܟ�8?��n��8�Ҙg��S��9�&��1��� 6��1s9B~���f�I�u0O�OW=�Kq@T���<S���R�z�K�W�G�k%�cŰ$q�pD�[k�q`GGE���}��#�N�]����&����m'���3��q��h��X2�1�����/�A�>���r"LO$ʕ�u�u����2T��+�ϩc� �!�
�ob-��蝄��OzD���ք�yT��/���!
�RN�,%w�,�)*#P��W�\Uf�8
 �3 g�l�a�	�5� ��AqMm�,l��T�tvҖ��D��.h��&�t��+2�x� >��i7�%ש#�=^�,���.a�k�I�>�F�܊�`L���ӏ��ɛ�]�)����#�a ?|��8=�zׯV� Hd5�뇖G��c0~��A.fUe����uڊ���B%���;ˣ"@f���D�����*�	�)��`A�0A��kn ���c价��|:	;>�>H��U]]���K�$�5�`E �B��7
��a�{v��i?�f.I=}K�R�yI�n%��_`�uoH�#���V斱~'Q��)Sm������>\�z!F.^'��\)0c��D��('��M9i�ϖ�X��jY�)���r!����~Rgfd�$v��0-�}5ԓ �{�љ���}hD�DB��`l�]��[�Q���q�6��s,M70,�)ᆶX�#��W�>��[s�>�{���3�Uru��d �hz�\&O��&����FD`
�{&N7k�k���c��ւ�Nj��}u��V��+�`,E-cy/;��O���M��5>��\�1�K�b���������;&��-���L�-vB���*^b�E�w�P���ƭ�Lrt��R
B�Y��Mu�;G���G]7맜` �=X�Z��Q�[��L�18��˥+]�^0�.��R�k�K�엎�����8"o���7�qs��zϐ��*�����E��2�:@���r���/yK�y/���&�[W���f>j�z�+�z"�z����-(���ynL,��L]��� u�T���XY�bK�3k���B_�ܳ��C'��~��x��T��;������A�ܾ�]�q*B�ڹXz�3Ұ��	��p��� ��� �N�O���T��cZB޶��1����%�x�'�").���� ��Ҝ�lWpcP//vNb���u"�ј�zf�/R�o�g�c�q%Z42��-���'�xifʹm���vH#��F~���zi-�S:������ø PeX���?��B��1��c�cʏ;��tj��N�b�i��_"�t<|h�_�V�!�F�SR��|�)O�@��y��B��Y��I���B���7�ۧ6����B.6��nێ�U��8��l@��\��"�=w_����zz�Vǐ5�����i&u�So%e"V���p���4�{4t/�����T����ԯ�B3.y녭ܖ��|��ἕؿ�d"�X ]��tu��F�'!\9�T��V��r��;nB�{���ܱy� �l}�ff��'��?�o,X:i<Û�j�6E������m;;eX��Ć�Q����j��j~���z|��-ը��g��Q		�V�摰�W/���NK1��w�C���JeuV�m��!��Jj�ʹѣ��~�����D�L��7�m���MTe�3�Ⱦ�aY�Q�7�C���C���TCC��7��9��-m<Z�E���%˴P�N�I(����MӔ͛��Ă�ց��&�w�l+Y����P�c���x�D�JL9X�e�.��T�=jH��T���B�@]ê���W3�1�	d�����������|A��7}/ݙnWIWL�|�(M�oyV��q3�I�{;=TK�-'������F0�:"k��L�廨V���D.!xl��`�o��6�;���(3ɲQ�Np0�>ѧ��9En�l�ki�ھ0�\��>�����h{���>�	:��n�l�|V����QNP��E��Q��h�)Л�"�SR=
=J�-��(#�W��y4�6�
a>�X�U���ܯ����9�daw��Ql�D#���w�ǿ�V_�j�[���6kVTb���ɯ3�����w?�+��r�g��Kv����թ��<_+%�ԝ[��g�p�>Z�1Rg�e��/�0�J'
"�@�������{�N��ߏW����Eԓ��`�gվ�^���y����˙�g[�:u᷈�b}n�D!���2D��F�W乩f�</��<Ao�J;n�Cd�@b�`+� ��"��)Ͻi�K���7��
�l�@����K�C˻�����O��s�E���:��m�!���_�:Ȓ+)�����pע%o[p�� ��8�2v�����?"i*.=
���g�3��\^r�فj���qH���֌׆�����E�¡��'�k(�A�2�Ml3s,w��T��C��������x�P�c���9:?;ڱ��(�p���s1Z��P�Dn�p���yHL'3x�%^FE_���cn�� ��
����w4��Q��[o��MR�� �9j��l���`�p��|���@������W�%	�̿�Og���.w�`�/�0�۟8�%%�v�y��v��5͔aK�"E]oJF�(�*K�@R3��;��\��'�GA#�L~��!�%�cpC�DC��ߡ7�V�'eh��c̠�yb�U���u�ԶG$CN.kQ�ÊΖ,���. �n���M�����ё=Q �#0.`j�$�18������H72��'JQ2�k@	Y������0%[��ׁN��H�@BuUR0s0�y�U6{�\Z��@C�<�6��Y[n�S�@-Ʋ��� ��c.\�=w8F�b�{r;�`_\Cv�m�ɿ��!+�Vl�!�*}\����--C�Q��Q�|u�X{� �Z$��7֎�ޥa��{�0�ŋ�?-G�*V���K5�����n���Zg��������p#6�
�{����,,��|_�#�!���f��ՙ��{�S|- }?��t��$��<8���d9:|u���a�*�b��'��E�����־Q$��1�EK�|{��:�Wv�C�P��|0�7��7���k�I�5�'��⦵�5�#��W���.{I�]:W��8�Ĳ8�eq4H��uh�=6N�v�=,F�R�d9�%���0�|�F���G
 �)ƫ��x��ѽ�ծ��W�OC�@rewS�TU��]��NO�N�X���Z�)����3Au���eUodMd�L�L����(�Δ�/~G�J.ϐous���� /\"h��*�1b�Q�UN��!_�����b�_�[;q	������n��o|r�d���4�pe6�����7U(*_9Kf�����:S��d��&*mn��1�c�AR�ѩ
�.�	4�u�P�<_�X�F>�t��b�[�C�N:���
�;�sno��%�;+#��M��g�<��xZ�Á�PxlM��!K��c-C�B����&A��Elq���Ts�6D�%O�`�~&�/Fg9�r�Z���@�\:.i�����&��}���e���tՙ}���er;4�C��1)Ϛ*GCQ�}P@��������av��j����E]]���.�F��u�n�6Q
�ט��@f�}��_���'ݤ1_��;hM��]D2$�5SL�u����m�]LT�����Q6��Οc`f�?"I�..	�W]�!5{��7��w>sqqb ��W��[�Kӣ�ͱ&K������mb��
Y��#���6�xC+H����=|��6.i��c!c9�����c����4d�p�������Tc���jAmA��`zq��m{U��c���kԜ�h�+c�s�b��<�O�QRn\ތ�F��_�3h���q�sO�i���(X���0i,��* ��n��y16��ި�5m�=eo�H�U�w��^��#���9ڗ|)cܕ��|���f����$#]��m��S��ǒ�|�(�Y�����YӠME�C�T��������M߽~A//�R�I9.d�{�r�$LA�M����M�
\���Z:�%.3��8M	���A�|I�}$1ȏ��Щ�(�R��|)��ؠm`q6��k�hv�j�.������8�&g���L@��=���QDʂ��7����5w^r,�)Ϣ�癓<��0�@#.󻭯�]�,��4�����=�^��`��:�(S�&S]Ƿ�
y$n�א���]췜�ܡa��h&L���nx~�%�k�����ƫaxǳm����w����1w���w������^�}���kZ��`��#;��?0���.M2G��M�שPS� ���[��"k��:ˏ�A&r�w �~wϸ�>|wd�Vь��a4dB��0�����?��Z�;�p.j���d�pթ��R>Ӽ@C�	�9%�S�[�^t�mN�4ÑDnؒ�������D��;>C�V	���E�{@ 5Kd���\z!/�Ę��Cm�-EG�&�E�L��6z��~L�)B]�)~�OQ}��y"��>�K}B,���:��bf!c�i�3W�|=����W:fH�!7�ˇ}�㦗��B9]������\q��5l9�ʬ.�6l JRZ�`ǿXC´Q��n�hͅm@�,���¤�c�n���ϩ&�6Q�����GW����j�U��N� 3t���N���j	d�q6[L}uz�~`w�^�O̹�|<}`���o��siB��&������w�rf7����������{cU�q)���+S-�xz����٫R\7�xն��dr$�R�e^3F4M�5 ē�H�_�Im���i���&c�b}d$��:�$�^E�9J<��������uQ� ��}�>���p�����7��/�J=:�#e��P�ŷ���>(��o
<�Ό�,�vPj@3I�dY��2B�wp�e�H�N�5ͥ=<Z�ׇ������N�0��I)J�z|�祦�h���Vm�l�D�u���Jˏ
Sw�­�7Uĸ�	=�A*�5ߪ�nA[G\;;v�ō)}"�KFx��p��UU��-��ل{�eۥG���:.�
�Kq��	`H�pA��9����7���c���~����F�+����UZߓV]�J���ڳS�K�������^�٨�9������&�g�b�l�9�h�wR���&S��P�?�doy�p���"�o���֪B��:k���g��������@�:�GSrNhL�z}�=O㢤Z�����IZ����0��[ǅ�X�\��^����M=-��zy�7��������'r��G7��^
D�)�3s��KG"��ث����^�ޘ��a��+�����J�.�f��d}���o
�M~�{��NQ_��g����}��.W�E)����ZT$�OU.�B��owͲ.��˝2T���y���#�%�GcȠ����$MOG�;�+r)8�=�Ǽ��j6w}���.�w�r#�O�� K�YX)��YY���H� E�����%���0/��j6w,EF�(E����*��7-����ⶥ�؀��?Ĵ��䏩�Qkl	�-�8bƧ�X�89�٦A �a޸q�5��ވ�u)��:S��K���?�V�ȫ~�`��hq,�_�к�X��<ۘټ�ٟ�k��Y��t��v�纳�X\L�l�c��)pr,n�ƨL�u��o��@��&��B}�`����hF�>�hw`4��M���P4!b�����$�>��>EQ�A���L���JӃ�D\i�_�W�>��]���P	:8���y�E���]���(�T[�r�h� ��~�+!�_%w��~�y���w��3Y�A�|c�J���X�]�QD<={ؑz��������NG2G�V��x�#�)t��ENL��,X��~���)����s����������~}�����w#�@��ѭ��H��׭K�'h���d/��EHD(j�r8�/��� ���ex4�X�|��<�zO�3�r���6M���f�W����,�Q��a� ��c^�� [vP:�����o@��h#'�nfN-�s���$����Q����X���G��ߵ�}�9e,zR��U0O��NIľ*���z�gP!�M�����P��[:�zI����m����((A����'G��p�DoKݍ�{K� �� Q�z`���;����_���k�f�Z���\:�������ړs�\���_&�[ͭ@nE-����$RC�X��i��BQP܅=���~b��97���DD�4�ޕ�䠀p��������u�	�KK�i��K�̄�v�G���3w�����F�n�(F�H@-�5oI�I��|%�1�����Ĩ�̻��(M��D�F�:^6�������^t���k���n�T�d
4^NI�2ut�7'�?N�<n*��;V9Z�B�X[��{��Ń��.c|��w��KN6}����07�d�Q�)3��$�x��D���E��ݏ�B���kL�D�!+b8c�}���3T��,��,�ڳ�"���$���L��\ҟJ�Y�1�+�]�o�_���$Cچ._?I	��ֶ][�F��{�9D'�xkh�߸����+�����rU��,�Eq�����*#41q2kOǮ;@�����P��.�� 1���h��γ������9�|[�x�(;1_K��`�s�Ά>��$ŵ~��MZ2B?�!~
uº��ې�T��zS���N^+]�q�Ln%��p��	���P��1�Db�0ʞ���<����FqRfv�'v}֞��h�I;X�7hH��$SKj��o���$��+�{BO�s�0�af�ڽ�&ӌ�Çǈ��_�(xݮ똀*�����E@?m�1��'�7��V��UL��\f~�X>����+�"���8)�o��^��ʻ	mqE�+�3�6Hd�j~]'(ЍPz��`�ag�2���W�������be�}ո(��'�l��-d�g����^�9���Q/���� I���-7��|��s=������暄Q_��i��b.�9���w�Ϡ!8C?�%U�t��rnx��a��s�&�>o�q��'o�ݯ�8=������w=I/��x�Ut�� ��ʛ)���e.$7��n�6�87�j@�l5$UT�-���gv7����>}D��>�?m>OTT+:�wͫ�y�k��Zb^�i<���@� ��є��K���ks�kˑ*t�owt��wܲ�ܕ0�W���˩��z�p�e.�K�ƣ����ǇFk2��STZ�9��0{g������������)�wv��Z̆������\��
�:o���=L��qv�w�Ҁ����E��S���Vo��_,'�B�韞"mƮ��;��&g�V ks��1yeՂ�>�ꒁ�G �J&��XLַK�T:�Mr.������$=-�&����A���a5��c��}�������?O�"�#
<ڒ�
{�5�2t/A}r��6Dv��4�nio3>~�Y�p"�~�/t�8��cS�_�k.2O�>w��#ݣ2�y�9bp�ܝ���J�J[5��+I3ɮ�b�����X.Aǻ�3y{��^+�HI`����(�UdI=3#�[c��l!(����h�� &w��F�݉���Y��ļ���<$��z��|%\s��=��v��|�	� ���3�+���b뷟��.�kP��D6F��Dq$�}6�����i������˽���?�r��$�\k;k\�gp��� ,F#ο&��C��y�b��h��c�dg[� 0bX����"{��:�w�S�&2xn�q��	1��c���O��}t2�V�M���ތm���D��Q*)�G��r�i^���v	�})���Bye�n��Lk��1��:��Y��iS[l�^�O�B�_X����m�dj��ǯN��]�{Z����y� M2�bbi����*/SS��U�mGe���� K4�I'�����ѯ*��G9dŶw�n��AOUV�㣞���7�@�����2�΀�-5�A��>8�<O33��wIq�����I�P"���7N~nQ�)���1�W�t��s�~G�DTÇ��u~��P��ͫD�t�_�z�~��:����wM"�\����k���̧������&(C�]�Lh��Pzns\3U�&G���w�A��V�K�@��%�ĕe ���D*H�mS�:݈���c;��!}AL~ ��v*��K�*,f�~d�ؗG�j"�ɹ���|���𽁧�*���\�M\J1/�v�Ĥ��B��"#UM�$~(Jx[���㈖����H��{� �</���ӝh�H����� �v�Q0�o]�"�=;�	��ǂ���s�0�s~w��qb�7�^fJ_�n�1�5W���4+%���$6q�4����!Y�e����yn�밼�h��r��J[iAK$�"��_��י�놥��W�ꫭ^��Jd�_#t»t�L�c�5bD�R ��:�K�S���?���Dz*��a�/꽝�b!�^J����c��zd�����q�V��4�J���m���!ٶ���\�-�KbU��qs��6����C�ӣ��!OWPq�}KѶ��~Y]�����J�2�����N�+8֕V.�yW���ܺ�U���o�yE�x��J��U��,�e�N�U�
��KF�����)Wkץ��2:'䷔�9����c|A�ـ���Cm�Y>���t���>3ץK!S����$G.��sY�qe/��Eńh˾�PL���w.�ڟ��N5�}�>�br�2���A��wr��e��+2S��sB�g�������7�R�*�yQө̓e�2m�����k�F�j�+V�L,k�1�U{�`&:9�\���Aj�e�i�����(;���I�ϛ�-�3�-�Q��8Zw�������q�	�wIt�Ӹ�'��8ٛ*�_5����~�0�y��n�����dM��8U���k���] ���G���~8���M/��M<%1�J��|G�^����)<��@���ļ1��9֞\���6����Ύ��~qv��#���F��d��a����<X���� ������o�7m���r����k�\R(��W�I<o|�Y��@_D�r m�_�U��:$O>�QGH쇢i�s)�A������2ʶj�r'|��V�5x|�y~���O1��j����t���q*�i�,g�Mw�/^���?&A�d"i=m�~���cK���4�0�,�x-��F6&��S,ңM�C1�yX��`Ê�r���̠�Ċ+�U*��p�v\y�(�u��h��1������1�'�l�e�mߥeoh��;�4ШS�f"�i� ?.-]��J�h`4n����~~`RH&)6��?l��]-@n3���noX��	G\g4]�+M���i���r�()�����ʷ�XmnAt� n[�I��7��UH�`ݺ}��k�����i��je��	����ը:._dDrjSF%�R<��sH�(�u{w'?�ea�~l\=��|-;h�aoŲz(t��o�wUHa�w����U0v�|0hl�S���~q�ӽ�jH�c~�)24�y��FF&�P6D��jC����y�y��g��74@������'��0c�%�/=���D�x�>HKŹ,/�0����z�+t�#U9�3�<O�mn��I� �6� �b[K�=U�-�#��ߌ���q�}([wj}� r'��������� �U�CB:4Ap�g颠��+��[�&���d�MU���Цf��R2�=�8��2��}(�ߓ��yF��M%D�+=/+�T�/��m'bci	Qx����Sn�䝐*<wBUz*c˖0�|��]IN���X-�u�j�`��I�ns��}H�.��e�/o�&[ �����3H�T��{�s�ia�8������#��i������v�g���6�m���\��˴6eMWeҠ���g��Si-Z��:�LO�,�?=��r���%O6z?�F~5�n{!��f1sc`@P��~A�f�ʺ��|���y�@���\��ǻ�=����Fp��i��W��mOd��$����*��r�ǤB>�7%G���ܔU��M ��Xl(�o�|eS��G���S�+ciQ�~����ڏ���4�򑪟<�A���+�Y(��k"�����dnd��m�a�ד���Em�?\�w�T1q8T�eXq��Ox���Ҳs"�bs.vx�4zg�����+�ؤ�:٣�F�U�<jh��Ѹ42�߼���22-l�Ŀ�p�`��0^��0����y�5-)pry����'=Í�e���5a��z�zǋ�\�1�u`��I�y%U���+�i1�<�	�pL��iJ�HS�uÅ�m.M��=m1������tW^�&������##��1�p�������>��M>��A�	u��cV��i��]qF\��Z�7�A2:�����z�h�*���r�I��
�q���:1�\���_dq��L��0�I8�V��#��ω)��o���#�۱���zOR�#�z}��3.�:J���q�R��L����~UJ��:ܫ��_ ��~&��h\�u�m��yǽm݅t�+�1��s�8{�~���p)Q�5�hK�\��%���F��ǿ��I����.��07���þ�4��uQ�����}*�<N3���'j�<b�`d�,��%�� ���F'�CZ3ԛ߭N\L�R!:�!�vD?� �|�ׇ�_+�����4�D^���;e��5�va����M~WV���Z�Uws��{��y}�X�/�n����2ht�kRSs�����*51���J
������&�r�̌��-����ڽ�U�u�X���Wց`�p=���(|��/�������U���S,� �z�v�^�C�.]�Ws�A�N�=/pw�N�哭o��e��;<"MOII�:�}�ո�5�gL�{���VӋ:��KxA���WE��)-ۊ�,��:�;o�΍/#�6���G��պ[n�}����:�I�J���bK4l�D|��Č�I[��v�k&N��#����5|	��!�J~gm:Uթ$���<��g�;�n�P��|��� ����'�x��n�[cC͜%���j�x��f)��oX��c�?]��[�wUanS\��?��>\�lb�졅�CU�W��y�*�����S�8!����"�>'����B3�M����|.=��uE�Z��yo�����7_d�������O�e`0n�\dj��)�9�G�x5̈́<��"�k�ղH����[��a_�Q5�y����ܧ�h���#����e>s&��􌚩B�ޮEL����oY0�}��_��E�_�4Ef\�X�C�!�^�l��ƒ�,�#�#o�.�L��9�ox=����k�|Z���K�o!�"��t���AY�}hY\������t{�y<��m��ѹ'򥌌u��z���H��ɹ����QU?{x71��=�M��*Fe*��(v�^�U��׺˜����#=�̼�޾+5я
	Y&8�4��vvv���3/N7��I��֦O�1�g^|w���3>��Zo�)�kzI�Ž���Dϵ���@���o&DH�?��x�����a�ӥc_'/�.�	�LF����9���1X�ePH!u��!Qe��O�<�Tt�n�dϦ>�!�c��Ox&��'����VG	�]�DB����*��ge=Ƶ������j �����&�0#R�#DgP����K�.f�9�9�в"�����MB��]����2�w�	J�?�p����Ak��6�����q��F`Vث�:lvɩ7�[�����}��#:��.$~:��I�2�o��݅IN��w�	Q�J�i��kE1�����"є�!����_$���5{]l_�x����*�kb�� n���*�12TDg2|������;��b�k�ͷ�L�'q~,̒���?�jM ��}��q������a�C���S��eY�˲i�ܲ�mP�;��'�22׉#��������w����~	E������@{NK
�?��L��Y���п��Y� �r���W�o�9�1�$8r���rV���G���eE~�I"V��_>M\��J��	�E-�RT8.N[�[��7����3�Q_VE�MwJw�HKII�HKww	l������n��ν)��s���|痗^��Y�^w�yFtO��v[^���P�1Ǆ������  _�(�q�cR�cyq�ª4��T�A�:��|Gp�~Fg0�5l�6�mk�o�!�e5�i�so*��DF�JV�!]`����	���7T�oX���ˈ�ͷ�����2�,cO���*���ш"�⧐Y�A�nB5V����~��P��b 3j�[�����t��n�x\��_��_6Z�36\��\LeW���w���m��A����0zB|��/% �,1�����ΰj�wh�F6�v�P���!���!�ˀ��)Y�C:]�CO�YUϔ�M��]j%�OBh˪�و�	#��pq��8[9;��ř�&Ab�ux#�)km��}���
��y�UŰ��O=Y��o�9B�����rc�%bz��{}��� �4�,{(p����;0�ΐ|�:�����g��$�|���E�,�=���� ��}��2�50����L�-ugג҄J���1w�~=\��k�G�_ȇ�f񵐜�_���RU�a>f�b� ":���R:�Ed��t:g)j@3�p�84xD-����< cG6
.p�a��`�eʽ��1�f�(H>�.}q9���j�o7Ռ�"yyj͑w��]S�Q��a�_1����f=��l����m�N%�D�PJ=�q����E��&3�4�g�*�+�><���!b_.+%Y�k��MK<�����򟕭�PɹdN�<�cֆ�1ux`u�����fJI��#�����.B7����b�eNB�<=g����˹������D^�_�&��'Ż�/��N`և�l\Λ5?^))�UH�m�Ӫ�g��ۼ��"p��ٝ�0���� �ي��V�c%��k�+<��{��Hh���+^�Ɵ���#9&���)�O�����\��q5q�Y���!�ˊ��&�}�F$;�|�<��ք;i�;��l	beb�h C����k	�R�ed�O��>��s d\�I�:R01�V4��x�u�Mc�H�Z��O�Vxo��xH2?~4�"+��t�a\�l�hs'����پ٧7OI����}��8m�\`v����_T��f�ۂ�_��T�({?&�N|hc$�P����E���w��n�]���;��4�12��#���K�� �Cc���=*2*��� ��C��Wk�4���y�.����g/H���U�R��t���u�`���͈�I_K���f�˫7��Zm*K~�%c�w�ʕ���)�d��.�P�C��v�"(�9�L�d���KAv���`�C�O��;�)"�{������+������^ѣp�vH[���(Ϩ�x8��w���^����, ���~�*�!��-X~t�#��*v�`/f���7]�����r5�����B� ���70>�[�ib�� ����W���?wGA�*ν_�����4"^�!X	���xP,;ii�}9�Q�K�G"���<�"�8��_�Q��z���#���t��vC�;IE4οȁ{p�W�ڮ��
/��]�w`�;�kP�uۼZ�EL��s�TJJ�6�Zf�˻��� �����rns,�c�Cv��F.���v���*�O��RZ�nVfQܗ����b��̈́�\<H��Ӏ�_8���p��x�H��()ZU.�*�|K��q)pA#&��݄�[A�����Ӡ�����I#_r2%$� �a��v�&nB�<�N�c��J��t���
���B������3�pM��g�)*��rKƀ{��"�_�������W�Iл�K;��̓i��!9�i{L'!��苰L�_~y�_��7���,��,�Oy;�ܫй�:�i�m�A��#T�w�:Ǻ+���v�>��a#WuѾ7ѱ��&4�w��`"�f6,&{%H���w�g�J��5?��62ҍy����!Ũ���6������u<Y��Z�����܌�)ˏ~oп]���"�:Q��K���uB��u!9r)-/��օ��&	�hi�[q� 3LsHM��[��u.N�@���7*�9��ی_�r�_O�1qU��ܵ��=�M[����ԛ�蹴�I���g�({cIT,�^D�W�m�M&���6c'Z�g�o#���@f��H)�]/-t
�����W�%�֨�4�a gɧ	N]�Z�C���_�2 �t�&X� D��{�6Z����w|a�T����:��(��
��`���䑰�ڛZ�^��[�C���"�f|$'�Bv#/�����C�-j�{u�b����K^CU���,=���p��J`1�&��ݪ?3O��݉��G{�qp+�6��C����Duh!V��/wef�ꂳ�J!I���̓��H:�rH2�3uM��`�9y�]��"����uv<w?�[0�s^E��I%�����;����7�������Q�ԔHLb�m1l�ƗQ�rX�%C�M�Q�{ 6���	�gvYn����A�3vif���1��4� R�;���\,�Z����Ã�>c�Z�y���`��b��3qӚ����c/3�x�������2<����'��Y���>NȲ�I�=/e;�&�\��ބ�.m���
�N�ǐ��ڳ�DK��[��b�������c���Rr�;Mx���_��FH�C���@^�u�X���P��#0�+B�ȰϸP����B���h�f�z<��]KM��1��׉�TjUŷc_D
PL-���o�/��E4�u��\��3SIk��h)1T��3�h�^�g��,�:+�Q"�/�y��s�5}]��MQ�!�H츢oͰ�x>�[zy�y�|�|e�6R�����9�$+U���o,=!�0K+�@��H��>Q�ZLI��l�B�1-�p%5;����H==��]�l^����;(!��?�r�PV���sʑ����� Z�$�[ݹ�$]�LK�u���	�ˈ}2F�h3e�*dp=�de�.�?�9;�9>�X$T��?(��3��j���fY]8,��Pq�'Y����m(b��U��tCCX㱂�1G"�{��i�\C[1�@l"Y�Ph'k�������*�X�Gx�v��B�a��D����?hE�V��������>AޒcE@�N'���sq�G����N�c:�e�Ea�g�h�d���Ȝ��@�u[n^���Bo�2(�AP�V\�?�~yG�G|y�g��b�#�=|0�"��4�>7Ǳ'�Z���0��[�88��w!�t�\���Y��il�)��1W�G�9����GZ�LSN���cY�o�3�_��|E&�-����t�x��}�`M����>Y��ꨩ=9�_�F�r��!�]0��B��;O��#}�0���=�������W�\h�o�?+[�-O��w['�
ē�:����掶m?�e��궎�l��SP���L���;��.ly<X�����ޏ�X'���qKmaF��Q���[�t��O7aC�(�_�������s��Rט��~�]NՏ�E�V���X���(l?�O�L�]'	q�� Ox4գu�s�������i5{�����������-%	�Im�����ne,[�e{����_r�U����,0����p����Ef�ؾ�v�?.s�\�k�v��˞f*z<�b��u���wq?�ۡ���"�c��8e"̣UcȎ��jF����L�Լ1�!;~�p�P��Z�y�I��+��Cf��u����%�qӶbx�r��s0L�*��Q�0�Vh@G����.{��o�Rq�fm�pY�b�L9e|�-c�%֥֨uz�����q����%?��_񻱜A�2����m�[A$�t
�G=I��%�� ����[�%1|J̌#$�p~>'�����f;�te
�%}�!����ɬ�[ǼqԻ,��*k��"�F]@�]'����e�u�ܘxo|}j��WI	-D	�*����K�R24��6�L��F��3�f�V�����9�T���;Sn���~w1
��dNЯ�H��P�u�iLe2v��3b����K���=���>* �@���Vh��(��J�0}���Y\�a����b��	M!��D�Ή��e��OUkʸ�GCuM�XՏn��zv�]���PR�Hj\�z�?j�ej����0m
Io^������_Hi���ތ^��$߁���q�:E�����h���d���9�G`n\�^HNk֪D�a���߄ѝ5��xI�$��mD�;ȴ�*3��2��������#k|�C2O}��P������B�I}��Y�H�Ã��{������kv������r����<�r���V�x�d�V�O�iW�'a_:m��bg�B���SZǆ.�i�1����X	=	�V;�G�����JR����c�A�/U�u�9-hic1v����K��ro���a�!'�vlY�t�P��n�8Fr��W���J[rfx�,n�L�I��穷�̼g���3�L熷�Ë}�Al&������@^z2_��Y���z�2�>��i\<G;���_L���X����P�u�q���J��R� ��nt&�UV9���}zA�K�w��I�YN$k,�VEbړ,
5�.��	�MU�5�VY&��+���W���C��IPg2:���Y���n��0A� �]��0֔F�:������w������v�{�oդb+��b�M��h��;�S�'Ba�wd�{Q�s;��җ4EH�;�ԈnAТy��YQ�<k�H�(�ͬ�ջ���K��Q���/Go*<]�?5ݖ.���m�д�5���֬�<�h2Jеp��(`�\����$\����cĎ������Ѣ>�h1T�[E�|cz���{ߒ�*ło���&C�<q�9[|��ۆ���3m?�v]~z�/�V����
��) c�q�b��X:��Hs�2u�P
8򯲍f�A�/�(�L��o�t@m���JW-4��5:�˳Ы��!?;�~ġ�)��u���o�CfNHg��J*���U�4=�hn�*�;�s؍����1�Ց��Stէ���!�p�E��� SC2��73&�7�����%�W���[�h��tx�ȏ�:/��ڰV��$?/����2�ͺcEk;�6"�V��V����d9�el��Q�j�Fۗ@O�G�x���C��UoկW#;'���_$3�agq��R^яz#l����� �b��9�;�>Ae
���E�Py�_p~���BBE��A��<�9�3�@�i�� U�j���/�C�Ͻ��~>��Rpk��b$/Es/=�]��Ӛ ���a���6ۥr�5W���Lu%�ҰG�`b^V�d�$�t�%�!�۹;�z��K��\�Pd�)��O��L�[^=�ߚ�u�1 z��0U�b�w~��Ӣ�C7�)"G	��;�t����^W�5�=Z|���C �d�3R`�����Ԭ(_��8�+�^�i�<�c���ՠiO���+LYC����|�7C^f�^�=jT�EL�5�뉳v�|Ym�^IxA꼯�k]�웟��u!ZĘȰ�/�����y3e���nl����w�zS�b�/��t��^;�{ć�Y����!I�=��	����~b�$�����G�2JJb�,B{��ǈ;����U ~j�j�]�����̼2�]�B?�[�y΃��*�ı�<��4qt�DWX������0�d�E���ԥ¿�΃A���2C����n�p�����Of8����=�ԣ����Nh��q�c������?�ڲ�C*]��czu�L���� �"���G�b�����\�����Q#��_�q���*s��tB�Z������4}/�qO�U�:`��t��K���KT�)�x=RDs�SR��MOGiq^p韢F�A��s��:t�6�"+�^א�2d�9��IFAMW��������^���Ns�R�Ϙ��ɆߟCF��,:O?��.�kV>�q/̔gL�0Lɋo�X��ݯ��8TXJ`�Ηۢ���0�'����"�*��R�GY۞:�y)H�y~��6͝H����Z��<���w23;��qI�D��zk>� 2B�H�$χ��'��1	�ώ�!S��k
��8�Ң��pI�UmZ0U�/�ó�����Z�P�T��,4kg5��v'��|E9�e�`#�7;��{�ԉ�������-6��4�����a�+T�?NIn�����ĭ�3�q�.�sb��2!�F��[!�\F�4���`�Zh-N�GJ�$��FڹA�
�*�I������,����a2U�d�����5�m�C�u�Я���h��&�����mT;w���σ�Uz۴{��WtB��M�g�D��"�X	�(~W,�0�R�� {�jj��[�-�w�uK�9���# �t�0�w2W�|A�Q(cr q��2Q�n-�w���MZ͙�t���=�0�*{�+E�t#y� ����M,��.k��(��S)
�*�-�|�T�:͟@������w���y���׈�*��Ą��02���!@�k�q,�4 ����l܁��G�k`�EA�=�u:�zh�ʏ�t))plgd[S��~�s�x��R�����#FcXc�;J�mz�x�b>�x�`<�<��fKA��=���5;S��O��%E� +�P�R W�x����7�t�bM<�g��HI�P�}��.Ow���i��#�<�N�����,3ۓ#wfJ�ߟ!?;"8$�[��y�7����s�
\%=�/�c�g���w>��[���=.�W�T%�f��o����k���y���&u�$���f���BouCBU}+.A���I
Ag�٫���w7T�}�dw�Em�Д�G��Q��b���D`�����-�S;oN�rzc\5���k�<
�E����TD��P�i�6�-GX��A箷0�=]��5��G����nǾ���s�)�VfMI^�@��9��q s���K@`��"�<���< �v��v���-k�#fB�5q6(c�)ST�3 � )�����;w�	��d����W�.d����=+�z�=l{���w�W�ZQ�����JէJ�mA'+�\Ŏ�Z�r�$�b���[���e:0�=m8�8�G��e<b�jH�hjv��9�sՋQ��L詛��B��L
�#2�.u��H؄�1�dމ��a|N��n���o�z�����:������:�:&���5o��aH�����済�a����f�� [l�P��$�B�VU�� ׆��왳�|���#��.U���Z̌X���Ti]���m�����yS��Ͷz�|��K��h��RtF����M�x�yj𸉵�yQ`����Ǥ��[����K<�f-O"4춡�֍�S<?8G��t.���R�v�NߛMOa�c=n";j�*1ߵ�_ב�Ep������l�ls�.�����|)"u�et�5���1�����Tȃ��c�Q3;E�X}�jb��r�8#ߙm��S���F1j^��X�ӳ��ݙ\%4�S�x��f�3������=��&�q����)�&��wP��,jȈv|0�bm����7���M�I%<�3}=v,p�bu�t�%0SXzx??���e����܀�`aI�U~$�g�Bd`Q��3��d��B�f�52VB�[�7���E�Ϻ'�gg��HB智'�:�I�*� w��^|�Uɧ���7��Ԑ�
P3��%>�x���.n�����%�8=�RӰC�i�֧�nTߦ��v\����eQ%�,��A��ۼ������6�<,:w9V�ƔA�SL1�q�ݘ:�������]v4�Z�A��tƐ����?˦��|�E����s��q�Z��S%VD���b�U��i	 �5L���솵K_��
Pj�+�E��E?7S�!s6Y�2�EՌ���G{��gq��`��v����
m�SO�>�+���f0濟c��Q�$�Gj��Q��'wE�A�bs��)}d-c�9��������V~�)�:�?M���_���ɽ{��.vj�k�����+E'��v˰!�-��P��kQ��{�vf/Z������r��v�퐕����uc:m���������R�G�H�^�@(N���>u�L���(01υ��g� J��� �:���2�`��L�3bV�u~�p���~0=z���~�
���q���/��ڙ�����3C3���i)˨��q��)�v�.�m��k���$;��nad)��K`*n^��W��	]=i"5�#�%5��tBL�����[�>?C��t)���N�ܱu�:p\8!�뽃bG���A��z�bL!����5��	��#BL������q� uN�r?	mS��}�������+Z��<�|��X�"c/�\�[tv��k�_q4�.�6��*{?�盎�W�^6���]T%M�T�j�7���EϢ8D�X�&�?���h���H��S����E�ʪ�b�O���/� F�S5�e��:i)�� v(i4n|�fU�z���g+�q�_dC��ʹ:<��]uj��O��yv�y^��X^����GV�TP�CنT�Rvv�W8�;Ky7e٣�,i��Ns���>Z�;l��r1]�V�%�2;1׎�}�H�cB2���@jF�p�q:g�����h���"�dR0W��� ����@���qW�t��o!*b��B@lk�ln�o��*�h���Qd�o�:{a�>Қ���v�:YG�?y�	n�U��f;B���֡/]���S�B��#�׋\#J��Z���O�8�}�c>�`6*��}�<���}�7�	-��k+�U�EF��*:�:�x�W�-$N� L����X2� ���bf�$����~�X��{@�¬M�{��&��=m������$�gL[D�9|r)Ƅ���y8���I�ky�pp��e<z���%Fd�j�m��e���<��Gc�u8�ۣm��.!=�sX���t�h$z�z�p�_6'^_�_�M�jw��p�v0�~�\tt�<2�ƞ98��- ��(�{��K�O3ae�~��O���$	rw�l�<�̟��a����j_ơwu{LI[ɾ"@x:=���0ۢ�����aİ�yA\�*l9��'ND~�d ��wB���J��z܌敳C���=��|ٻ��c�2R��ۋu����� W��MC�B���͖h[�Q�Lj7w�K���u�Sc��r.)��İ�+o��o�\�U�fe=.M���ĕ�Rn��E\�'�E���V�l�-��,�G�ad� %�����ڗ;�<4��MQ5F��uk#���s�f�]pE��X��8|9M��F���%��	9��3~{���'�y����ov�t��)��$F��x Æ����G����8ɩq^�g#���TṠ�wZ����#$F�����k�&��.^���Y7�T3�?S#[b/2�PHpU/χ�T����^��w�,��n������fW����h�V�/�X	�$du���L�#�Z��������<�+��^*%S 㒳;ܥ�?��g�w�rc���a'�Q~y�{x~�.'�g�A]t!��vo\[Ll�~` �X7�W���P;�9b�3ܲ���D�׹�k��KI���I؊䇏�W��'���Y�vﺔ��kk��b�Y[���o�@J�q�NOo�&'��#Q5��,�d%`�����Ά��a�r����x����H�Z��WP���˱o��:�������8��2�>��R�s����.��a��ȏ9�z"��w7���c�pr�slnEC{,�v^4^൚�6܆������P�*�T�zZ�r���	%��x��2 _2�#s�4�>t&3�9m"�o�G�l���R�'R-�6�?�V|M^�[�N��=��Ĉp�����ŶJf�c�]PvD��������{P(�k�p�a��G.L%�����'g/�����T��c��0jgTbm�Ɓ��`�֕���B�t�ñCڒ,�	k�Uu�o�r�s����9^L�C���ls97��u!�V�1ܽ�a�������N8~ �����dgY�A/����*׾Q������\7��[�������o���^y"d@U+�u�n` �4|�'���7↳�:�ȝ�m���C����bN�$���x�{q)%�ut�C�\%w�3��5&����� b�+��~~g+!�Ϣ�NǸ%�Fυ������$Kh%�����I��*�N�3��Gw~0��i���{��ޒ:����cJ��2wMQ�o��gm��3���8m�����jhI����5�(ѿ�ې[[�2o�Av
8�O�K��H�y������*:	jFL^;j^��M�L������6XR��Y�)8/�z��2�7Z�j��E���V�P����q�q�o;�8�9�bB�phD�][
B^�/zʅY 1��H���<�������w
s���ڬ(]��v��9�s�U����{^�<*�(E�Jw�5���P��\6��l%�JX�Ov6�?`VC�?�<��=�J�&��x�=����l����Z��~q��u>��3����_�'K��qW+s$�H����L�*C�n��]R�IS�=���7W�"J�Y�n������������ykX�Ձ��l,��ݥ{�����T���#��ˉ�'�K���>����,����Z�	EzЭ2���UN4��mO�)�z�)S����q�!��f�#��R�d�Q�QE�RC�R̀�"��۫K�$�������k�~��-�:nwT�j�]���o��`<:R�Ʒ�0�Ȳ�^��QS捿���<ɋ��(h"NW0���9Oz$�~���Mj����ʏ!�1/'W�N�,- )z>S���ag8���� ǹ����L�~��i�SDH;�s��[��������â�\�q���z�Vv���C2T�/�����EZJDN������ab�7�P|h�.1�(���y���eI`�N:Q
c�¤D�p�QJ�7���L1u
 ��o�nl��PuG�nw����݆{��q	�����{�O��:?]k��⽚�ad�U�K�x�c�9�,x��hb)�VF��=�h��@,Rc��b�\���$��S)��C��d-"TB���*��WL�|�����1"T?o�xW��b]?�o�ܵ��7}�o�4�/�Q��%W_�iQf?�۔���2��T2�;RX���6X}uB]�O��z$��@W�i��T����]�~��7~����G`4�d�xY�1Y�|<,�X� �LTR�p��ǧg1�0m�� �����B{���ڈjO�����U%��������r�qh��qƊج��L��/56��V,.�"_M!�k�
ӹY�t��\
�=a�f�EQ���\����^ӑ���3źc��߮��b�N�w�Y	�n'��i��	�a�!"ȏp��v1�ϊh��R�I{w��{��=���kޚY�*h����g_�W��I8����C1%��C
���N��ԅ�i��:V᪈^���U�[I�bMk1�{b��9���+�Od&s�7u��&�@D��7������fM��*UA�wj�mC�(��4�����e��ͱ[u�;�Q��{5��d�k�k�K4]!7����f��z!yޱ�=�`]��n��e�|�d��]�Δޮ}�`�.[r.l!�d�|"�ј?�Y�������{T�Dmȓ-3�����\o��!0����������t�Vc�?\'qR#_�����@Ax7��[q��m��ք!�E��Ds!���s|�3�_���l�B�G�����۔�c�q�?��P�P:��p#����)���Z�R��u�C�5���k+aB6�^-M�|{<���љ�o�T����Ժ0+�:�2�T���E�B�A���
��W�@�%�؂��h���aZ;���	��`�'I�@#���(+��:+��� ��dX�?�,��.����ĸl��*k��������)��\�����g�\��~�6�	x�1GG���F�-`~?О����C�H0�ih}gH���G�sp�D�=�YS���bIp\>�~ia�)��:���{���5��+�یꂆJ׵C"EH�t��<ګ�Ӊ�;���tj�Y2�.G���_x�Ż}��p}?��[�ŭ��ƖO%�U����}Q�o$��q��]s�$c��񾥙P�����`|j�pRB��6l���7;;JziO�|)�N�x<�*Z�~B��,�����?W�>�i|���A�=� ��<�/�j��hu�dO8s��hZ-���[�̈���(�l���u�_���z����e�C�HI'O *��q����<���{��[a�� u�`�]m�x<�
MOKi�߁#�ۃqI|Aq�5��'�VY��%c9?'�ؐ�N!-x���-�Lރa�Q ���1G�>��pJzf�V�'Pg�N�����1����!II]8�{r^�N��u����D�d�;��إ��O)���HzZ���p3����Y|�zZw��:�uom���"��5�����#s)�F��x����˫�2���	X#���
�G��R�P��=�W5�o�yl&�(�֊��.�u��i{zD�O�33��,a��4�O�/!*���2�T�`��bh5x���3�B.
��P�:�VD�l� �8�5�8��uU�}�j-��y�u�'�%�t:i?�b�����Ӑ��ԋ��� �p��}lcnX^ԣl?o�|�0J��[��k�#���d���T���g�Ms�G��P>�� ޫ���Ȋ�hܱ57��K�y�0� �<���a�>�R���2���S]O��U�W!��Nfꢷ���cr�DK��C/�	!�4�tm�1�L�ٜ�*�lf�����H�`�S�$z>�9p^T���`s'	\��Jzt�B6r�sג&7�7v�D�K�q�c�â1#.�b�v�l�M��9�zk)�����=�y��x��.���Ś	-��]��"w�9T�o ��[n����	%��k撖]����&�N���ER�;��`�ܠ�C���e���Xn�@:����L��{���Xǰm�CV�-USf!�Ս�<�LI ���z8E�h
v<�~+���#0��PB��on�N����!�6�M�T����
���HhȨ���OGF��g��o���`��L�`!h ���<۰���(W���.-�V���k��g���MŔ�#zmL?*���1eE�����w��n؍y3�c�#�5��F(��Q��{:f�m��\����9|��j���`"v�b�c�w&M}ǐ��cB��^���M0���˲2&J[�ǎ>��N��^�h%meN�0��|w��L�..� :�F�<��kB6lu���8��Q������JG*�xo5պ�����~��hԀ�"32.^�JC8J��;����DE�G�c��7���c��*^��O!�.#a�f�z ��9=HϒS�"�m�P:�_9�'���i�*a�v���]�8�8OG�d�3�����m)<j��PF�G��y�3~9���6+��G��/�~^��W�3f_Z��E ?��2�o%x��*�-jtf<�����ד����11�?���	��0ՏN�	�|�8��b{��7����j��,p�t ��~�쏴�{2��t�3[Z��:W#ܕ$���BM�%9�x��G�bFg��`%m���,](�Y�Q�.��G[1(*:�\�Q�Jh����<|��էnUM��Az��޶*D���3��k�	�G�v"�A`�88�0��%9;���%��2v�I���	E�(h�
;Wʭ�ޭ�=����窽<P�� F��K��$ԒU��P|��Y�۹�<ہ6ꌔ{��]��.s�y����7om�$�'��!��?�-��1��Nxj�<�?��;��<����������blÉr��u���l������in��5����w!F�W�|��B�e���
��-s���(��/��n팸���iX��߉?����^���D�6\�8~�����F��kz�.����{U�S�]���ȱ�"�qHo���F�q�R��X��$�Sn+�O9�i�俸M6��:����dIN�F�ϗ�����ahRq;�T��/U�q�˧�R�\�@f�b>��Բ��0��;�6"���6Z��A�I�N���M�>�6%wLO��
��<�듘�FKg�K���ޒ���c�����yX��96$��\�⍵.)1d�0�ކ��Na6�XK��o��?��� ��f��/r�$6&d��mW���Al��f(.���$��f�%Zo�t���-�������[OZ�aȄ�$���=@I
�/�t�+�{��l��0^�-J^���b�Y�I������S��z�zN�����۫v�Tr{
��#��j�w&%�e�ǍE
�]��l��l�D��R_Gpeh��b�4'�l{g�ۻX�v{qg�L<1��E�$}�9�r+b��mÐ�B�At2NW��e���w����ov#=ڴmd�/Z�Y�C��rKu*�����6�Br�HD>6�}@#�,�@��$�"ncX׵��f����,N��Q�4{$�<$�|�9�J?���ߗ��w����,	��rc��#�*�"n1ѧ͓Zu�R0ԡ���_�Ϣ�V���������Y^���`��pm���볞�F�R�(�6���
wm���Sz��ڔPن�*��A��dI9��r�s��xb�OIA�(o(z�H����^�+H�O��΍�,�V�/w�����n^�%?�<iѦ?D���;���
�� ��"�d=��1��>�h٭?��S}O
�!�"�"o��1�����I̞L����R�ҫ����#���1;�]�M��I>)��ww��0>�NÂ_)���j+���}�7���C��Pg���mZ?����W|�����e�ֳ�iB������@����	r�ſ��y���A@�l�>{�%��l����q�Y۞E�CU+"���������b�mwW��S꒓B5�<G�yp�y���4����/��	sW�"���֤��9�ȫ]4��}���x�J�ϋC?� S��M?i�(F,N�/�(<�n�E�|b]����=�9z�}/L&�d�\�6I�wk��ßTX�9��w��q�I͛~�5�D)��u��햩���p͏��_��q^����O�z����Hh�?��-�}�H�N��Jnŧ��p���%���c@ؼ+���9�t]�qt���o���=*���A�h;E��̩I�W�٪�+��6W@�DH�(8��� Bo����!685�뛈!����n�B�D�~r�^���$t��g�C�:U$�A(�BN�M�7��Z%0���|k��,�"ế�� �M��z�)��#�53&I��~�.`����F�V��]x��#k1t��,���Ǝ�:[N�̀@�
���� �_�Ǖ��ޮZ��l���WV����ȕ�Ƹ:�tW�H��LS��H�>%<
ս1M���+%���L)$R�N>���Q|wv��F!j�#���.*c>U>�H����|�>Q��������ד1���;�4���dXe��}�,���W���i���Û��t<^��(4�}�ͦ�5����U�
L���?<KҌk���mU���_Ja��E{�B�.���|7�G���&�q��/���M{������T잣-O�X�����.��:b�<HSi}���JI"��7j�B���]=�8O�gy4-�u@m���������TT��kw-��na2��Rُ{o�����g?f� �:�������|�����C���ͮ����⋃���xg�'�U�R[e��'������	]ʴ�ۡ�h�=X���9�x�%*eBx�"y�l�Kt�n���,⭾�-����|����a<�b&���Dz�\(��h�����ͺ����F;���������`�g�;���1e��,��O|���_��Y�Rx ZMV��b\R��@9}#_I�i�s��r��t�F3�0������iv�M��c{9z��{�4��Rմ���|*q�u��k����	��������q���"q;�xC�t��i�6#S�E����G�LG�?�5���T��S�:�z�=�RH��#L��s�my_=K�S�O��OrB��9�k0�����)#��~�M�w�#1�t{J=�b���>���Թ����ψ���"�È�7����⡧���ЫD��Ye�*�z�u�/���9�й/��Z}0�1�����%]>��|ݲ���g�y$Gj}��%����<q7N�p��A�'*?f��ɚw8��6�?{"ąR�"�	�x�_cI0���9��1��رv�:[G�>5�=G�3����)�D�a�G�_���=�jIvP}(N��p����k3�|�~v�A�$�2�_�-O!FZ(u��J�ʭ>�+��|-.��t��[G�-�D�Z.�e�
��B�X�T5��&ƣv7b�&��wu韯4BUMkF�⃁�e�Eu���?��}!&Y�َVc|�)A�8�����y7���ӟݽ%�yh�~���l��B8Ƈ\����O"���_��l����izݚ���o�B�-`��,ԥ�	���D.)��`q쳓��Z���[�
��k�̌/W�<|��<�g����3s��I������?�p�5M<����ӳˌ�h��$�k�*��B�5�t�;j �t����(�8QMHٖc�n��FT���j��'K]ͳ�ɜ�D��`_q��5��ɘ��brz��^gs���-�B�wsz鵘9� �s�g2Ӓ�-�pl�1Ȍ��b<�aq����y�d�}�����5�t��@Ѥ�ԝ;?��;7�:z��A^��ʬZO}�ǔ���[�`�4�uTT���A�nDB:�K�N��n���SJP���������}�֬5�uO���ϳϙ#����?b�I"WX�{?
q��x^�"X��_b'k8�mKݢ$n��,�?R:��q���g��Lr�Q�����wZ5;SbL�z8?k�my�f~����>��P���iZ���!��W_�z�ߗ�j��kw�-���k)��`M���O���ѧ�W�n�k���_N��K�R�7`�j���w��tK��}�B:�ZR
w��k�?��G����3A$��ʀ�k�}�xT�IǮ��|6��(8j��/���췓�w>�!*V����\W�sF��q/�7P9���c��\��X�`o�%L��}��q�:p�Ij�����@�
��526X[�]²�D���T��/�
��mw�쬐`�����PO*ʭ��r�0 �z���ן�������t[�\T0el�=�W�b��rZͪB�}6��_Y�N����/􋱀������bB�F���)H#{��f�l�)��&b��U�+�1�&��͐��:�t���NZ��c�f32G;>d��d�T+2�A��R�ń�UzU0˻�f�(�+S����t��?W趐��|�j�����Ϩ,+�P��
�zG��k�c�I�ђkk-�]$&�S���}Tmt b5L�`�%D���Ԣ�1�K=�r��nQ���e����P� ����(ք�)e��N��ʄ?+����1d��޼��$���
=�����A?k�?��� N��a��l�����}wji�Ƥ�*���_��i^܃gv�>ӧ��kQ��;I���Wt��%����~��BDsl��X�AY�:=��h���ؒj��LՍ��;��.3/��>�������n�V��06�J>�.����w2!- �6@;8jz��BFybuBT��
��<��LYc`��
��_c�G��D��j�3����b��z��!��B�k)�T�>J�#?���������X��ܐ�D�	��V������o���1�n���-�z�1��
T�{E�@C�GX^��d��*�o���%E���ղ/I?t��p1�wѣ�:�&�2��a�\˘W|C�8hc�&���Χ]�ؼ���-T�'�wz|gp�|�m>���o��l/�r�z;9c���H��l�2���"�zo/����� �<���,p��9����aҩq�0hh��`�q�O�%�q��-�&��So�(��ƻ����D�.���7к
�}��խݜ�c@y����5��2l�ߒ�0!�m嶩͙���0lq���a��o.�G�c t��[�[�ո���K�WT�aB���j!�k
�������1���u�5��#�^�:�C-C[T ��k�f���SN��n@�[��)aNO9W�G����/j��Xq ���dn]���4V�-�ѿl4������j9t��o�[�)�$=ɝ��B&�^��&�%���!��*�s+8l�/(�h�"��ߍ��ľ u�,T����l���O�e�L��@�QIY��LT*��,�a-���pin����N{;�]�k}g
�Nϰ.�K�Z�'��T�[p;c�z�/sQ���}Đ���O��+5H�ޞof�ݶ�ߎ���� ��uΒ�3�x���%;,�1{j�}%ʓ�|�����u��z�u�2�8X�B��g�x�|���\[A���c����]����TnS�BwE��P�QOp�����>�vf�mI+e����~�A�@{� ����.?=M;ag��^j%���$&��}k��]B3�|��c��{	��K�/b���e��=���K��'�������g5�s$6`�*�-s��䎿�0`>����K�S陏����a��@5���~U���ǋW����(k������JM�UE�cJ�WGX}R4ѶW��Rȵ�/+!U�N�Qt�V��R�k�]v3I#&��0�(Ɛ6\�`��$�#+{	�ʟѱ��v�Ap����և5/���Q�f{�z�B�Q���s��Q�oOt}��a�i	/S�[���d��L�B�Ξ�>��� ��n	^(�ٹ}X�w@�LZ�Թ�!0�2mh#��,�Dx��x.�5�G��u4�?F�}��7�Gg�A�&�c���?��ܰ)��ҁ�y�CL$���1YV�p1A�<�Xwض�[sn���)N���kT��Lq�i���Lgs���S�e�3���#��pB��`�(yc�ɳa��������g��m��+�5��gO���}դ6��n�?��/`�ɍG���_3o�F[n<.� �����pP�z<W�3�Ϧ��WZ*�/��/���I�׳����:�U'�Ya�Q�6�4��D&�!��r�v 5�=t��8ȸ��ҙdj�]��YfO���/W����_(�*RJ�?�?뮂!�*!��l�ϡًA�٬�?��"�-���#�Pl-Z�?��gOe�c.�P�/��9�R8�G���:>��k���E����կ�~{n{&���^w��d���	-������h��cKp�`���"S´�5������^�0�8ǐX���_�s�;wZ�{����Dn�� �5'���uH�%�n��
&������|�=KoaH�s��wm���xVa�<Y���z��_���a�� �zRsoE`g@�EY�[֘x�!�%[�):��Q!>�r����*s֎��P��$��L%`2�ZZZcˋ�N��0O#Wo�E��ҝ����'%�r�c�HQ��w��=X���Ɩ���F��h��W;fg�
�E]�\��d~f7?��Jl�ŗ��"x��k5�R��ސ��4�g޵z�dܵ�)!�䧭�57��Y߁�x�$!�F�=�X�G���^��?�D���6<�zV��ݓ�<���A�s;��o���/V��A���
zּ���D�|��EW�K��jp��(ʳ'j9f??�����ދ�@�Uso��h9ɦ��&���4U����f���� ;vzJi�m����i3AhS����=�.")�s�].��ݮ/��~ka>M���1y:�Yv�K�-�<���JvuFc8Z_�0��_�����S: 峪�==S<�-S��_8^54�y�E0��_�q�����xo�|�� ����C^�"!O�B�\���� f��_��r\�m��毱H]b!S�����I�� +W7���0޽iu��[/��$0UL̛�J�S��;�nC��֎4�L��8��%�V�~�$;�S�L>0�$�f�q&�_RG^�y�Xs��!&r7[]K2i>��(L$z�@�4R�V���W=+�|t�>W:4,{|�a;r[Tձ{��&hʤ���"�`ǲ�jZbV�<��#:y~[ő���C�uh���(�ϞSay��n9+(>f��v0���PU/	_�q�Zv�t-ݷ`���Hjַ��A���t��1^��=!S�A�}���Ї�u��sfBg�?���N[X-����G��[K�d�2VuTښ7Z=��UKDh���S�	�&�є�#�e�h���f�**��ֆMǐ�+Nf&����*�,'��=��W�qP�8�=�0U�]���Bi����邼���1��u
_(5WL�Z���W�=�G���_8R��G�hԎ�}{RQ�e�'���j�9|�Ie�"����M��T�>��Ȉ�nt���k�W�������m�3r���q�v#fˣ�x�~r,�ʁ7s�������j�IϽ ���1����sΦ7�����X�m�֕�=�I�
)@�3X#�}���������h3~��IJ��ð5c�l�u�fM�s,�͵{�,��?"�G�$y��������q��{R��1U��?w�^c�na�9��oQ�ܼӓ^<-��A�:{��3u��"(�����]�c۟�NV�!���@1YQ���'�/1�:7���^_7�%n��i]��B'k�`]h'C���y��̵�_��sJ�W�2;bT�緱�+�Us~S��R�]���Q��T�����|.N��(U�qӣ��L�}_��u9�!
[�w�i2¦Q�Wgl�NuL��c_:b�>i�����+�X���� /�5Ơ��(����jغ�4�G��<e>kiz���t��G9�(�ik�\��-c\�N��Δ��3�)��M�P09�v�+%������6�6���V�'-Q��#Lc1�Ǫ)}��2�Fqp��X�a#��dP�����ߢ�qV�/�둵F��z\[��1L�D���z|����\3��<ˆ�����/{��s��6n�� ���F%K	�J�d�ww?6WUPG���x��v���`��a�7������Ƕ�Y�>����:y�a
I��z��h�3��=9O��`OD���b���7Qt�˜7�~/�������͟x|����X>^�z�'��M����X��7'�#�p;f���A��}?۽M�c�\Ow[rʩ���ӡ�%�����pi<����k�9r��-���X��3�q ;��`		>�n:�E�\��Vm�!�;zJb��:�4/��h���HB������:]��H�p�,��$'8|�k��Ѫ�>XO�
�g��!NL��O���T/�Ԋ>�x�5�Y���؆}�ɞ�Y ]J~��\�$͘��!Jja�����!�������jM8�Zv g|�"���˻w @�V!;9��n����+����WoD����eb�a.�;W��`R��b��&6�E&G��.}�dl�S�w��OJy���
"c�*��"Av��2ƐhJC�_�T�BxU���L�ܖ��c�z�z�6W���3��p�ZStX��ia��8�y��e����=[0w=S��@V��֙�#��H�M�����b�X���nm3���{>�����;��$I���LT�!?G_F+��.�3u;�e���xz��5z�_��Q3J\At�WK�r�r.d�$��݌l&�9�A��0�dw=�=���0��.�V:@d;���^ �^�=3�QF;eI��L%��19�2�~�4���}<�m��kl�z`׸�	vWB(S	v��	_�h��]��?\�����.KQI6����؀è<����O�E�0b��8�@-�0�`g%.-VV&������E�|��H�j�ſ���8�+8BŊ<S�m�|I.�GBj	��x�^b�X,c#��d�������q��i��XB�3���ґ�Tڒ�"�*	�l�h|�*aҷ�V�(J��t&պ�l!׬F7&�SrW:��k؊k���Ik�:��izc�-�d�v�$��5�&��&4�#��֪|t����m8�`?}�c� ���$gb�c���)gr���ni���u	�e�:+���ԏj9ʕy��%�u�$l��G��" ~	 2@V�,Fm�����_�H�����Iip/�FB�3���WT���B�N��	�rt��|��z�]��8�<��z�N���w��b����&���1���h�e�$OZ�i2R��I�Xݓ�=L!�߁�F:>�2�@����. {T:4�%n�pǟ�U%V�>��%�
[�}�X���k,!*}sK���6����J߈f�	2$m(��^���6��ru�(�������D(���w����=8"oD��{w{J��E�a\n!ar`n���ê*&0gSΔl e���u��f��rt(�M�\j�v3�G3�U7/M8�J��Lګ|]�NM�G�Z��p�#/��Ȁz*�*�$�B����G:P�YI��}���~�g�j�O��O�)��#���X`���))��_ڼ r�^>��Ǝ�F�8�,���2 �;���X}ڿq��7�_�����:D��Z�Նǵ	۬��$���%e8��e�]�C<���Ŏ��EF9�H����\@3�8��-�� H�H�%+�P��U�y�+�֘?~�m��b�GE� K2�W ��/�}r4F�I?Ԙ��Z3杋���B��Z��#��_EX��
�#��K��2�_���u�E	ڙ���)�5�b����U���F�;��q��.-���>2���EwRٯ�fk�܍PV3�1:��ĳ��W��4v�D�XZ/�B�y�=|6�*����c�x(�ch�"~�dXEP�1��#� K��h�!�
|���"�o�F�/a��Y����R4ʗ`!�x͌�v>��=]�`�{qU�0q�~:Y��6rC��L@|%��CT*�d�J��4��h���V.wNⷶ]sL�%�>Y�4�1�F龷�0�k�8��
v_���v���)M��c0G9��,M���z<����!��Ƿ�1����#'����ſE��W�~�	�8fW����#ᘄ�s��g~�Ur�LN/��w���-j&�h�5�g׌۵љ�U��K�J�q8��N��z�0N�zm��s�A�O��¼��n@6yi��N&�_��-Q������Ԗ�����!�<7ĸ�������-��Ѣ�joW9i0��gP%��;�-$�%��$�O�-V��LJ��!Y?�c�Q$�S�N��.�Z'+"��B��7�ĳ7�<�vo�ޙA,����7�ٽ�!�k�>+ǔ�!���+"5��(�}��|��.�\�
q���B�v��=�
9��m���8f|W��mҳ3��&�.��&�*�ܲa�7sY�jč4~��7�Y>f�M��?V	�3��F$-��ZFBoKh8����
�z�����E^ֵ��:��������s�v!�!n�H�Q� +�_��
s+��'r#��'��@�]'��N���<R���M��_���^gn���x�R4z�qV:��u���}hTB��_!v���u�=��ׁZn]�"
���L�+�s�G��4*�[�`Ǯ��O$=�ô��Y5���q7*��Ԁ�0_����d�?�8�'���1s֢MB�ڢ�����Z�:���M�MXSU�x����C��[�A�w�AՖ#%
(��2kfW�kb9��&q��k�T�&{v��'�������GV�'|H��T4�'�~L�j�ǝ�ϴE�Fd-6�"�� £֙������"S���_�(%AYXP;�à�T@1�+��
���ʌ:�����04��OZh9*�!���◸B�����ҷ�a����*jѳ��y}�g��OS�ld3V�s�����hغ�&�cO��_��%+쩣�"0��(�"���������=�f�ͤ��	V����D������Ŗ����J�f�{o!2�N�6!Ϻ�(�4�Mf"�e�$Π[�<����۔�5���e�ɗ��]���p`8a>���3̓��\lQ)$�����؇ݪ�Y��*��2�#Ľ�{ӧ�*;r{c��'�K/��f&�C��mC�$�
�p(����a�^@�Q_����$��޸����F�d����p������L�C$�'8:���b�H��$Ҕ�[�<��F�ăC�ZG�\p�--�y+ͅ�{u�D0ML�Ch*Ʀ+s��(�q��,(o�����c.�U�ҝ������_����6Y�1SԨ�?�B��]�(|���?��J��&Wqfh��}je� [^�1C�����ʊ��1;RHm��1�V�*����/���ݲ��zk�Mn~=�7i��JC1#��F�0�f�ey�x����� ���DRAm��Z�Ee��2ytTĦ��-=�GY�s�J���&�B��a��8v���SC����b��!�&L,�=C�͙�Prz�*��:�)f�7aq�r[��]��B�=If�6�7n��%�:���h7Mޱ�����:��P�M�]���y��իΓ�����݁?��\����YO���y��b����ą)�^[>� �g�⑪K{������B��$,��-$���'u��+GJ�e�ޟ���+!Tb�>%~�=-��|�{�a=�U͘8�y>�k�F%6��VN��6C|l÷W��X	�7'�NCX_G6�v� �2!�������ISH~�<\� L��g쓋���#�\����$���n�#n�{Ug�pH�T �-�j9�᢯���-MbhT4H�"L���e���:�y:�.�H�g֯��o����;��z$A�h`tx��wTHɗ�s����gt	/���j�粻��xѢ��b�%F]r���g4�7��
UG�1t�AkI�I'&p��D�4���"���$!&m2��y�pb�I$�IИ�����|٤�����$�Qٽ��Vxm���{�H��►$�0P:`w_�����9�6��kV
9��c���*\@��j�9yTɞ�^ϛO�zH�����Yf�Y�9f�qG�Q&M�O>���UOw/9���u����bN>��^\QQ��������׎-�@}tѠ�ץȚ����")��w��W�B��'��fK��W���4�ΫPğ
u ��/?���;���sX{:�;�rE��	E��PfM?.����cKᖾȾ�0������<7f�(�g�<��퍳�pu���Uo��q�(�'=�����.*Znu�4������U�=4]����8�x*h�Z��.!w�{�K�M*!AEF����8��t�S<�W�<��Q?!n��Fɑ��%���J"�/�&A� w2�Q~�ͭvh#^{��jE)Q���&A���Y/�(s����cG
��s���V��cz�X�&*�߬Jp���fs2�	7ǩ��U16j�0p�������2�:�F�bxcv4	3��!�f�sƚ,f���=�(P(�F��'��ŎK:7��ev�����ę�.J%���hL�q����	�E\�ۇ�O�N�"ǹp��Z��vN.b���Hp���c� g$;y�%�z�9�~R�$LNկJ-ʠ���g�L��[3MG۳r��_���+-��55-D���Σr�[�]��#Bɯ��֓1���w��T�VUn�l\��1�~�]��a=\c�tӚ���/ҀtH܄�g�S@}�.A�nw�J{[o\�r��8�sѰ�s�DLq����Ҩ�~�	����J��K���̳$�4����f�?F�1��e�,=�r��ZV������8���r�z9���=:�'%��f��`�� �#"��0��d�F�_��]��|THEj���gN���j����Q�1=8���e�^���Kp�Y�����?(�>o3��U�e�U��v�l$V�9�B<�X��BZVy�d�x�3��&D���BOZ�E���`&�w�'��;��MtMg�{V����|����P�+=#��zO��Z�(H��?H���}N���@�H���=_��+�(K�~
�ήb�������x�J4?P5g'��]c���{O��h��E���yjȍ�~W�|VT
��2����==�4NE��,������?|po�5G�����xI(����	�<:�~%���cˈ8�'����'�.�:b������p�����0��,� ��u]<¡�n	�������bN������R�<�a�6�y�oT����̩(��&'g��G]���m]����;�4��\��&��ݞ#���HC[���R��1�T8JJ��ZR�l�����:ė��ke�gB������-�;{_Rɂ<0��*\�ҿ�ф�0U�Tӭ�KE��٭��[��Ċ�w.������vme�q��/b��ͥG�s�^fi�� ?`^����5�J��V=b����ޗT�0�k���H4��rR��Wg��ْm��U�Yb�eBN��I�0B���m�֘�~'��:�Z:����ZL������,ٕ��ɽ�3�qp
J���f��Am8a=��-JZ5`�3ĬA�a�^�K#٧�[pz����)����.�����D�Ԛ`�����x��av�:_ � `3�-}����R������2�Z��r$�{���8dkԡ(M��w��]+b�P�G�A+��؅��A��}L��Ј���}�i8H?���	i�8�^�],�t�y�oR�_4_n�7����<�y�~[زRu$3�v��g�e��|{��vB\����WbckB�x�w�۾�������m��v�+s�&���L����}!��׉�g�s��b�(���mE�:e����js@R�r�ϴ�؈��Z�U��E���?��g�0�O_U���z���� :GB�֊:���t���Ϡ�����h�tl&.��Q7�G���K��a#���~�~�_fQ��w��P�1j���@H��520z�ʅ|� �g5�1�?��R~�oS*H�ޮ�~�����T�3h��@�Sw2-�M���/���;Uv,�ގb�LqУ�g��p����h��k���凝�vL/Y)&~��0d�hK�D��ߺe��d"S�ǙZ�T��A�w`�)��*��u�U\Ds\��Bu�����A*A�mi�(�~�Y�b?��D�x)T�._�����/�j��d�#Q֖��%���C��|�������z�SV�`���@�����E.�bF�%X(��M�+;G�i���Ew�
Z�iw�P�=���yh7/��}��|ڽG{��RkJy��n�hs���-�+�ytSCS��o�.��P"'[����/αDnT���wI�,Ii���;�Y��c���q�x"�l=08O�Z�RF��5�s��pC�&w����"D��A<�C����{~y�#��{ϖMxg⚀�;�E���5J�-��&'~��2Ct��j�T}�\���2�U�|3쌍UpKS�}�冀�y�?���kc-sP��
�@�h#
��ǥޅ2�SZ≔�X營�7�{3�
�} cK{l�d��%��3��+����"v-�}U g��n�|���3TϪ�(���@e�����ژB��a��L�:A,��nijz����i��t����i�r�y�h�K�\�������{.��ԏ-.�xӿ�O��D��.��9P���Z�]��Tf�#6���lT_�-�	9*�����)����G�o(��QM)�<P�U#V�U��N�nj�;EL�0�S*����G��&�9Ku��V�xq�:�z�;��n�nj�{���>:��B������?δ>Z�
��-�d��q��d*x��h���1�Y�����ɯ���r� �ITr�)�������橍�s
*�N�f��p�Ƴ{�	7����waʎ)�Z]�7[u���D,��iw{Y�z�08aOS�gx�#��C�n�~T=��u%�pm%�y�s��*9��둽�;���y���a0�_Ls1P[�@�^�����<�8K�qn��a� w��p�*���&�f������'=�n��:؏�_-T��leH�X&'!|i���)kB�y>��W7XX3�3~���4g��e%��Yh2%� �k5~�C�
�D|{�pZ`�XX��ީ}�`��Q����{�j�>Ţp7��n���Rj0��]�B��Ytv���o��n�&���7��8t)�P�Lb1�dʩk=���G>bl&������ �Y�h���j���*�(�?5I��Y�*�0f�����k�K�i�FG��r�а�y� ��~[dD��1�R�,W��*��Q�-�c�_:I���j�_,�!�^d�"X'�Xh�2��mH �J���Oy�8�w_GA:��g��C��n��������i��2d���;��i���Е�h��av��s��)��G~�k5Z,��hc���D�y�_j]�[�}���r�����a���qrW:����G���$G����2��rg&���d��GD�ؿ�:�7�=	[ܶ��lh��`�{�s�WTu��Ns���a *w�f,C��tt�2x\f�������ɻo�NxF������P���R?�W'������l�t���_?�zڤc�z�nn7bw����V7%��'��I+��
���s��b�tn�o'ߍ�$f!��]Ӷ�^06!R���~�4a?U���p�(��A�9�ҷe@���b�;� :;��X���g�5�4��U������FG���0�_����G���[`'���k�l��x~X	���x(n\�x��r\#���t���m��gD&��<�/����Eu��Iϩ�ʶ�w��AȢ�p�bK��.��˦a=B����{@�@��f}��*v�O���V�>e�١T\��0�'.��㇍�$�k�b��R�y�<5�:"|�繴�6���	h^
rk^t�\������0'�`����J`��֥r�Vgo!�<^�@�b�5�#]?�h��`FG���$�4ʅ�ya����[�`��&ݧ��K3}�i�Z�=$.�vk�rX��l1�p7�E9��j!^���An��}����������O��6�����O�9^�j?�G"v�'㹷�j���
j}�����Hy@O���Ul3Fa�*���ԏ�4\��j �>��I> h��B|�*G�g��Z��ǯɦ��~�د/o΀���6v��4*ʱ��0�*��e��9p� �O���[�:�wd�v�/��9���p�F��C{ŇeOއ�g%׷c<i=P#d���W9\--�8bJ�h~�7�����B0��2���;��8?\�v�s�B�k�K�r�&ղ4��t�Kg�qs�dd�I���p�@Q�F���Vr�R�/5�����'6A�`-��Pnc�5Dqㆅ�۳wK)�9W~j���;bR<�1�E
�q�!e�Q��_G�Q�
�bn���i��>�4�2AT� �wi$�_���ה����u�^�5�*|�o����ͮA��G2��I���1��U��H̩ �6й�^`�7�4��|#�#4�f֕��;є�~����zfOLo��V�G�P���E���M�O�4�*��_0F-���r�e3Ԩ�c�Nwء�6�T�/��h�Ώ�qn\<���OU�oP�[lS  &�u�|R�1����Q�A��p�O���}�����;ja�y�T!@W�ZJ�؄����������*�.�	��3�����.[v/*���2'5ͯ��U��G�i��K^=�NK;��=����#����MU�B=�TX��w��.h2��K?��{��u�yQ"�gc�u5羼�|R�m��D[���d�mZ5��j�FfH�q�͐�$��Y7��~8�d�U��� ����Z�w3�����ehb��c��>�,�x�)��<*/�������U_�ٸ��|�ܕ<���>������<ZN'o�S	L���%ơ��'u�|Ӧ�/���|-h��7X�QU���P���W�!�5��h�j?���+�����ˠ����:ʉ}.:RŖ;f�;�NX������J�]����>����kk����O��|K8ۅ���ľb�s�u�?b��/�I �!<�k����:���1E�&�C�^Bv��c��ٜ���� ��
�9\�6�ۺ���jZɿ����|'�*�׻Y1R��$�a��S��l&3Gn�TLm�P���on�+�p$=!����k$�P���f%�H����Ya��_�q�S��+��������,6/�4'k 6'Y�����v���b`Kg��%*氖^���}�O�N,{���Q��r#��d�XMq��_n0}���o =s�}3�� �.�H���j^gf8��z�^T|S��(�"�PAZ|a��]�Q�bǫ�-��VZv��!#��|�2���~j�壗?E�i���IMO���oIӖ�������=\�콟A�8Z�؅S¡���]:j|r"-�����Z�G�1��G8$�L�3�aPJ�O崚��� �տ�W�<������e�2'v&����eZB��K��7kX���)�;8���1]�p�\70��CDQ�{� "�N�&B��~�*|BN�1��Vߙh1��R"��p��3���.�2������k�M�m��gY�����c?���d�ɒ��ۛ#w��U���{��u�� ���/9�'�'�D.d�A3$��y�33�]�U���'$���c٬+��ƾ�5���;��jg�������<G-��D�u
�W�s
Xw=hƨ!��1����n@�{�(�;�nz�%���m�c-:��
�J�̩���ų/���'�6�1m1mv=aZ_neJ�(�p��u[��s�A�����ܛ��k��JޖLZ��������E8s@�_i���������W�&�j�'�z�es�$$x��3Epo�P��{z��?:d���2x��H�w<�=I�J��᯸>��.1�
�����=�Ս�20Y����@����-�93�]�>|�wl��(?�9x�_Kx�ZL������� @��z�G6���;>q�������lVL�]����'�akg�ac?�`M8^)��X�s�2��+E�α �	��*;����FN��L�/��Xzb�����Pb�j��	s��.a�=)9����l|�Uo&�4*̐~*������@���H9.���p%����� o<{�	K�7{EFj�A�Gex���s�l�z{���Lr�����n���^dt�K��h`��x5P���
p����y�t�F�њ���*pz��)M|�Gp�%��oH�A%?{�|�O�����U��^������lR���HA�D���v�ʅ���2�Y�� �d�oơY@!"Mo�'$��:�m'sn��晩��3܇���a9���܊��$ߎ�b�?��j+�ݻ���<~���8��#�<Y�}`���ޟ��J��%J�&�PWb���is�x� e��7�\�G<��pw�)�諴vT��7�D�f�~�N�^��5�I"�׊���k���A������:�("���<��⻅�%��gKܮLB�"�]���n��}���TH��ro��X6��N��+���k<vi�C��w5�K��/��ŨQ;��Z�h���RO���K�k�Pz����k	ţ?�ΥS��_`FL}ry#�wm�/���`gB�-�zSB���GEFA���ނJ��C^���S=LGBv����t��"�\�T�G��>�_X�LŐ�v`@ZsAv^���2�f�ȸj�Q��[M�/o�e!eh�F'���5�=|���E�#y�?� &%9{'3Xŗh$31�"���t�����I���V&'�_9�X�>&�v?��Nr5]�JHK�ћ��o� �X�R������44N�X�Œ�JG����
�y���Y4���4��`X�5��i�u�(d;�����ө�ޏ�
�`�%B�->�����К6E��6i�S�g�&�d�ɖ%�w)����+J���%d�2	�~(���D-nM�N�G^�I	G^|s/���k��<b���S�W�����6������.�S�ɘh���#kED�٭b�*��U_w^7f� ���w���s»9Y�،��yt ���񘸴n	,�v�ŽC����ڊ���L$S*��A�-|�AS^F+�$�(�8���J�����;��	E~�Yҽ�G����(���UZ��$;�al���6���Vf�A����9��uL��^@RQ��F�,�Z�T!G�zfԲ�w9{c��xGA^���"R��N9b摚�9��3<w����?$�>*,��MmĿL��#�x�&���8B\R���wǁ�Z��^��o^=؉���f������ ��PVX��w���:��H~��5�I*�p�BW~
�on�C�9)�Em�A�5�#�7d������<v�D�Ņ�{wS ���2�,���$̯\-�s�Q>{�j���	�65� ����ݞ�U�b�z�%�ԋG!�.�)���&Y����,3��%���q���WA*x��4�5�ߚ�c~����S�^��$5���y����8�_yi"X:�D����jmy�`t��<�� ��������D���J�h}���g[�tt��次����{�����hoO��&�O`>y�#�^wd\{/l���z"�ܿ��|'�$��]X�Dzg8�7�
�L\g#�I��I�?����a7J1[�C����qB�[�i���:�"��C��ۿŲ���ǫ��J�F�iEVх�ȶ�r�,d �8��7}+�/�?j��g���}�h(����F�����T�;�0�����[=`�
�V�f�����՛̀U�~�D��9��U�(#;S���U����7��f6�2�Qb���8��p�C};(r,Y&��àB$B�1��ǹ�*�#�e=^����#B�3�&������,\u^>V�k#X��i����Y���r��)���P_����"��q���{�Q�0}2P�p�n�PI�����Y�[���7��:�T����1�25�T(�K$P��LG�lvR�6V;�K+�wpd��J�S*Nh푺��u�/sG���-g�Qe��^�a=Y��n{1k:d7���B&U�יDl�u�]�agR�o�������J�F��w^F������о�{Um	UUzN��-��w�a�)�"|������|P�B��렦�C�X��èn�ݒ)��R^��*]mIm~Ҡ]2k��Zl�=�@HB8�����5���w��~���V�o�8W�: �k���Rr��+�}���u���?K}�"Zb��	H��E#a�>W(�<�G\��E���8ʅp��7��%�+j&�᥊8b�TA�n���ǂ.i4"���$vn��$�9��3j��$�j�� �����cTV��^`e^���	�TZ-�5O�v��^,� �d��zпS���W4
�aɮ����I�m����Ys�mf�����Zp�p����70���9e8D+E���P���{�F���ڭ��������ҝJH#-�1��Ԉ��Hw*�� ]
H��P#HK���������k���s���U�̰�z/���t�n�gk#��uN���42�r��/��.⓵��6�fmzpS9:MzA�Xzw��>o�M������ÿFs��!�Wl4mX>�:_��>3p��RL���O�$�N� �L����*`��ϳT�k�[W������?3�2Hտ�?�:hO�<!���'�+&�1�����i͢}�~�����?�]��Oj�"L�'��n���I�#TF���Fλ&��&��,�K�,5�86��Ԕ��W�������3+�N��I�K�6$J7u5�����|I��M�M�/X����J���Ki��ފ��t��+�*�{�ʧ��)� B0,[M��+��)��dGjS�����Ε����!�H���!��eJҮ9��2���, s\wMf��Z� ZulJ�:�U;>�b�	yrH���1�����b�������Om��e�gbC;ɕ���U,�z���_U�� ��W�T�zk+�ڒ�%_7��J$\E ����\�VOoln�폒3��p�{^����PῘ�?�o⮆�{������[ޗ��UYJX��	���1�Ǥ��<�?ǰ�ݱ�1?�Q#Hr2�={�de�9^n��}ȘO����o��ј���ENd������  ]�)�Y���d#s�w�f=4���IwѴ��=3�U'e��>� �2�^k��R4K���׸�yrX�V��\I	����s.�JB���ES���_�H���堬���%|q�����௻���-��#��j<��c
	T[L���{ytүցD�S�SK)TVVYҳ��l��:���r�� B�I� �>Th����GP�U�at�Л$Uދߏ=NT
�:�Z,�����9gՙ�x ����9u�3��W{�~�T�n��ܤ9��r�㒶Y{�&x�M�D3Ң�w������7Ci��!�r��|u���[�p�`��2�k����1�͆�}�J���u�o-n�Q��=������5�Q�c�&��âaʍ�A��W|�c?�V֞���h�Gy�J�o�
��-��-��2:�|.��5� Co����ɮR:A��n���VP�i��'i�c�U�0��3-8f`�Μ��������A�~j���\��Ol[�����Ã�r��*��V9Ĉ{#�|�Qӊ0{�c3z�gI�F�RTx�X����B! ��M��B3��=���y�N��X��B��ڥp�"��5���UrC���N�����$�T.ɼ�S!@5}�o�O����ȏ�+���q$#�.1��n*�o���n��j���n������{)�0TZ~�����8Z�8�7��ԄV���Wr{O?j�����Pʒ�a�O���R>�q�UՑ�[�t�=�q��jA�uğ���񈩤du2���#���mq�����q ��`Xi�B�J�!�ָ�]C����nD��݂�3��M�\���o��(Ꞝ����IF�Ŕ�ͪ�����C�q,1��_�j�z"	�X1��T�9���%�|���qY�䴢�-���]����&]�M�f�e��2N'k4	���]�d�5�Ì�+
j�p�5�/X{�=�~��c�� [�e9y��/��lcH�G�`��~��C�orz�7��7�$�|��5b���M�=" ��S��_�9+�uřl�8+;4�߯b�ˤ�St}�����RFh��Lެ��@ʸ���L��m�y�
�3�����vK�v]�����or�^��B��P��^�A��o==𗧙-(���U��eC�U�1T��6�,${�f���7��0�W��]7��D��	��h�t�I�T�{���Yj\4�܄ ��y�d9ɜe6���#��3�ϯ�G��>)J���ƁUqv2ӕ�[���+s˰Ʉ䲽O;����͍��~B"z5.���-���͕�.�L�;���Y�!0~x����R? |?�����C�d؎۹���$�`U��'ߚ�WI��N�B��[�h�ݲ���}����s���񰬦�k���b���8PR6�x�8��K���o��׿���j�
�|�5�;�{z�'�\�M�<_�[�9Nm/V�gH��8�6�:�0"�]v���+�eN��]�/9�#1��V��{~�C��0r�6�����'���&��!�t��Ρǌ[����گ��zۙ��ۍ�RX�qq���>�=���^⇋�ʗ��U�G�~U	y�<���<���"�]:I�tL�q��T���h� ��.��9���Uf�ܽ���3�1z��h|*J����A�����`bSg%�E��>�L�6�#e:?�f��j����`���F<~�06�i��(f/���I�N�u����rױ͈xq��|��bGj!�W�2�;��3���q��/�r0�z���{ԻO��w����Ǯu�5���@��w��w�
"g���i!�j��Z��� 9�ǲ��b�w��U������x��/%���mp�Ͳ�5�UP��#���b��QvM �Ro�w�!�����'ZI�1������+��T�����H@h���g/���>xo��=}�.���^��ә�O�]��G�Y��[�+���C�dU<����?������L��Ļܣ7�z�w��s�Uc����s p��;��pqw��[HW��%��Wle>��S4����'�"��cqXct渍�[�����?9�*�)�T�T�%�I���&�	��h��d�_���P5�-�R�}e8���Ɖ��i���Ѳ��2�_���p�x<��1����б�c���1���l��J����e͵��j���FH㒃����c�c<zpL47�"u@��dK��:8w�X)Z?sC��%����[}�Ux�/ЬK�d�&���WA��V�5�f�P:M���b�U�؁����a�%�T���	�֏5�!��ޅ� ������V���QW
Zt� �z>%K�*��KM`H���4}mQ:�G-�<6z����E�����B�^ ���&vL|�#:5�E�
�����H祬~�k{\�8D�������ȹ����J�� E7B�5���ݤq(ŝ$���hZ���*	3+v��7��eo���s����kRj��D~�vv�@�������^���c��CtD*T3�F�f{�\���'�Y���j�L�&���^�:u%�DOX��lV����-��r�K2��)zX��C�=Q�IA^�]�8k�_��o��R�����S���b���u[;��;s/P����>�&.��M��a)t��:��VT��I�0�����C��v�b�R�ΩO.��}_���s��7v���-Q�m��GU�E���h���Z-Ԟ�^���С�C�dH��Q
s�R��If)v�(w$�UD��b��5�������R��3��6�: p��nh���`}�!�&y7 ���z��gEG�b�I(2���Kw��"�$Ci����N�7���@�R�Ą ^�E}2T:�,k]�N��iWh;N�假��wy�vת�Uu��c�YvF��V���L���:��a}�Ы��g�{7���%&�f��t(�gOW_�m��e֭��_ͧ�DG_q�m�}t�Nj"H�*=.����� �^�q:"G�
T���#Ǯj����?;�N�mߓI�HzB�j����@�K�߹9"#"ش��(X���X���9� �z߀���4v�ѣЫL,p77��`�����?r���sѹ�}˧����0���J�ZϻH��3����1�b2y�}z1�R�d���(�$�L��t���L5"l'�O,h���kv��N�C/���R(B�.����fdl�D���1��{5[����ϧ��7�ϩ.�n����2i�W�� �P�y���4����?(���Vf��<AMt���t~w�EC��{���{OV[� i������fSZ�t �C�uJ��'�x1Z2�"6�G�^Ll�9��\�=�"Q��_ Zl�)oγV�!���7?�r��o�Xg ����QE;ĸE$(�D����P���ٸ;B;E�u�76\Ep�?袱��|��-�#C��Uo�H雭��n�r�j�}D��S�^�?���g���x�D+��h�i�d��;q���w�4B%s0h|
�녴ih��+�g��[��k|�Hy-
�z8ݪ���Qp8�����qY�,�#D�YWp	�az�>�=��%E1�@%���4_�}?;CA(�	���D�^ 1\S�~D�X��>�Zh0[96M�sE��k��}G��9xjO�@�h�h�(���m]��C�� IX�����a��| G�����}��T�?V�-�]b���>Я�J:(c/D����	/G��m�GR۪�u1�mL�m~{��Y���7��Ol��]�L�����������+�+��t$���VV�X��Y?!���5���Iq��10 ��n ��&�'m$.�Xɛ�t��&8�m��`��W��F��p<�3?h,��Z �&�����w�?���=��W�q��hV��Z�����z���P�=�0�B������.�q�9!,O�g�'��ҿu,��w��ܓ�p���m������ν�����Ddp�Mзi������Ď��ў�5��m����3�H��,�>��<��v�Ā���?�N���2��Tθ%R�{^�ƅf,�}1+�F���vC�_�v�&h���]/�[{�O��k*8�O�'���P!]�K�/�_E�Ur�h�<0�X�w�hr`BmA���Q����dc����]�����oB?tC((2�r��R�U�剛�I�>[5�+�L�u���K����� ;�| Շ�ָ�!y���Xm�Vڊ:#���ņ�o=0ó:�0��������R�+���20�)4�Sl��>��y�����_��S��qWϻF�e�����<ߠd�۠r@<��ܤ=�*"�B�>%���/�����.
RWz��\��W���D4�q�'�_�I`5JӍ�A��c�S�hD0�j�:����	IU�'C�����������2dO�����ʫ��8����� >[DM��4���S����R.�/����%���{��D��_E9���{�!���KQ�"@���l&|��>��*���#�|s�m����l�&�/�)�[��D.G��^~���1,� 38��-	��z ��;s�;2���?ֶ������IK�&��k����*s�L�ۃԖ���{�M�D�<6�X�E鳶��F_$�-��f&Qb�:"�\�$���4�C�>��_P���<��k�6s�ۿ��] i�c��!C��#��BU�`Gf)�<�T� ��J&�A�/ԣ��a�vn�[[���6��A۽M���٭��Uc�\������:J_��a?�`K��s�Uǝ�d,�A�8�� D���=��ޠG��֒*ϰt�4�QVc!ޣ%�>����˳�Ľ�U[|�C��mP8�3�DJ���_�a.wY��U{s5�ى���Fg�Mh��K�ů薙Ď��������0�wwXz�&=�8#)�֋�P}�z1Y.������3Z�3����u��e��ahv�x�u�*\��5�	 H�^�E�α{$��|��L�6��27���}�B9�:C�;����0v~�� ڹ#��s�����iR�:/K��7(��8�5���:.���Rn����,���fCy��g'� �o�|Чk �_��&]b>N������@�U#/�rq�Gu�hz��!���e{��������y���s�}�s�C_<�G9`�1������څ��3ϰ���v7�u'�<�ۼV;��R� 9j�yam�U���(NK ��F*��u�k�'"5�����>H[%�4���k�Q�tK"���u+�ܥt�>cN��SD���bod��z���I���򿚋�u�S�U�����`�'3>ay��<�5;�t0�c�}3ed=5��D�\{���$�S ��C�]��͖��T���)�C�ܠ�ո�JjT�Y2��t廘�}g���s��vTr���-z8���FX��%&��(";f)o�\"`U#{o38B5�l��x���|,�6��ɅPr��{}œ����4fW��%D�t�K��*������)�%��clԕ�)�ܳ�k7��#%M���ɹ��1͕ϩUfe���̿ iQ�Qm)eҽ��N4�#I�e��:�������؝�(<Ә�Sk���T���W�N�� �Z*��y	�a��Z|{�s$	״��������~�c�����gr�`"�.���n�N]���{�2���1��/��Q�m��0½����W�Q�@��:����b6��P��:�����ה���`H�4`���!MIM��r��	o䠬^,cP��X ���
-aW[�]5��U���[��̋���,�fhR�M�����aBcr
��
!x�d�_h{t��fL���A{.brAe�bwVcX�im���)�9Hua�:���`g=8�ux��`�����W�x@Fć�D��PА_��O��
12����O�^,h��>4�p�h�W��O^j����x��<��J,��]�S�n����ƩUO�LBI�� %ƛЫ��Wi�SS��J�eG�n��VA)W�9��1���"U��Z�֧ � *���������,L��3w/��N������z����w��L�2"�|M�@��3����w����ߎL%�P��&z�`B#�Y䠂cZ-��nf��v%��o����:�J����Y0�V ��>S�hp1Fm��0K�g�i���R�<��#z�Z&�!�d��ON�l�9��rXug �R ��D�g�E%�a���I"1 ����c�A��+zzU���-��/����3T���#�!p����A�M+#R�9HUuߏ�s}x��B��uCOY�� 07�����H�k�>��j[j�3������2����&��?�� 7�\fٻ�pK��;��v?$�Y*FXQC���l)�A��.Ju�¦�����=�88z٤<��0�o'A�	��
:Np�eU.�as`m_�#�(�ώ���<�֖'�?��M]�=}�)	�e2�u�nf��%�9���;2��T�?����/�8���n�եr�N�p� �;�ޚ&#Tŭ� _-*�����b��?����E�l��ŝ<⇬�"Rd˓���x@fY�q=�qM*���d���G�)A�'��wS[zn��b�Zmx��q�lչ2��$l�[@��j�ɟ��������쮽'�H-���3Iw�=��3�>������[ܿT��`A��}�߿T�������Bŏ�(��8��J��ly���l��ͪ����nc�r���MI��,��&E*V�}}��d�t$��e��Op��z�v(�?Դ��Od��e��&v�e/W�j��E3{�7��i,��یo���ވ��8�
�G�
B]}/mݠ2L��"1������e���}�� ��c׃���np�^�>Y���v�	� Itƭ�DW�ͽ���0������k���]��GH��sw�
��O��X�#�6�m7ƊƤ�� ��~�u3�6���.����ڊ��Iș��st&��]�r"G-�7s��Il�8��GP���C�R�����V� X������>B0��t��� ���{#���>Z�e� ���
UƬq��Us�B�;p��ngCUZ��7���M�͢nΒ�	#3L�I��E����}C��`'��$�AD?��o�m49�:|��$����-J�)�#j'�����K���2Lz�&�i�҅�����i_{�b�5Y,n����J
P�:j���N{S��w;&�ߌ�;��d��g��9u��AԖ2E>K���{�o]V<G���59��6�^�b�ς���oz�A�;�c�ݛ��`�����I4p����U[������б���F�I��ĩ�z~��8�IO�ȃ�� %�i�A74�4�8���U��S�K�D�:��*�Z)Զ��꜉�(���6��GC��ȃ�6��1N^]
�ɺ}gkJ�I�b�J�����_�2[3~/F�L����?��}Ȯ�Z/L�J���:�� =���%"�R�g:x�vo;a(�0�EV�����+��X�ƾ�\�6�J$����dTN�ױ!�*�ު���s^�Ao�mp& �/���q~0�FR��{<�KK�w���{" ��$!(g�?-��Eed/��K����:#S'���X�~0�aG��_�*�޵B�[)��&h��Sɣ-��|���~c1��WtRO�ŏ�4��.=�x3��h�Y�L�s��R(�;��4Z傜�t@S�o�2?̞�����c��j�&�?�HA
C�%����*�������k��HB[�ڋt��iu*�X0-y�7�"�8z�.߽��Ҟ�R��)+��*���v�z��G��:S�(��@�m)��ݴ ��Qy�Nq�ƾ���?\K���˜�=�<�A2gT6���'BpJ��W��U�{���8-Ҟ�:���`�ޥ:�q�� Zf�|~�h�SzuG�F��?`��op��LR�
DQ�5.=~�	��.�]2����m��ы4U�9���&v���MN	�DԪ a�2����)�u~�V Vϧ�V�na�234�c��+�?���[NV<������q��	�u1���;�\f�Ǉ�ql	��
T3��uM-py���}i�������U���<���W����e�n�iH���"[�L4��"1�!��t�q@tqo�#���ӡ\j�W�X!4�-ߞj��?��ǦK��*�l�7(}�[l-�]��cZ�PlDn#�6�w��n�}��k��s+��}5��t���J�[?5�*@��~g8���/{�r�X$]n��s*s�<�Z����:*��l��^����Q%P#�d�o���oM��H{�d2��4��7�32Iy� D�A�v�9�T|��'P��kn���H}:�c�_� 6D�Tt�L�M]w�	'��m�[��۾3֥��اa��sp!M��x�oc
"|nK E����7:����SO��c�����YH��7�������b\YW��!e��~2��(�>�_r��W�e��W�޻9뽦Y�1�&r�g"���X�M$d���w���ݸFDY%�Y���Ц���^�	��ҩ|4���bڜ%i]�۟�?����<��]˃b{﷍h�3Ko�(��2�Թ���)e�F�2��d���Ǥ3Fe+��z!��c��Ƿb�x��13�\45AZ�9��S{Y��K��i��}ѶuZO�7�'�PP�t�3!����Sk_'�(<ݱʚS}y'�Y{�&�1�1����R�C�FqV�qyv�_�B�X�,{|E��ӎ�o�v����#�A5� J�L�Z-Ļ���%JB��Z�.*6&��þ�R��`C5\|�>���5WƬݮ��f)^��R:��?N @�x�o�-HM|�����嬞t̙�S�o��E��DVA�<} �;J�%r���ݤ�.�C��^˜CQ� wL�e8a@���#�9�ɳR���)?�W�$l�B��c������v�i1k���*�Myˤɪ�_�K�v����ٔ�B�A�Y�gM�߰^!S�2V9X����?n��*`�j![��S��g�1O/�kT���� R\�B�C����Sw!���۵/�ȅ��f2�)@�%��sj���~���W���g�sJ�?�/�2�✭�F����nIjm�z�$�h���_ �_��?
���V����YЗ�ZZ�b�^/[sn��κů����}	���e����2��XK���=��B�k�~K���F�b�|B�ѫ&�LjrV�b�(��Ζ;����'�����1��^��T���%1z���-�fF��
��ߪ=ӄ��6&�슈�)�{���ࣛ��Aea�ڤ���P}�ǫk��*�F�x�l�KyF�ߙ?���EnY�no�SפNy�$1 �57�җ�}kȴ�����`�>H�`
i����Y=�#5x��k��Cg�L�i�q�`�����q��9�|���}��f�����6���-�yAc�[��P�	�^����}� {����"������@`�1Xlb*nǏ��������U����a���	��;H��������5A�-|�NtoiN�#'̼�y�B"�5�%�|��׼��:�z��}�����O��#_��"��!�}<zz�1�#��.o!�%mk���(�9���}ɤuA�H7dGg�}h���g�Ak-14�����X;y^jV����FgD����T�������~}Y7��iU�|'�իM��`�	SK-F��.��K���y�[�w4����pu<;{��T��i�P�?�R�Ѽy��sצ}�m�#"`���^(�p��$�yS�.��yy)�->2D���
�g�
N48��l�'��;��|���o�_8��TѸd�o����2��V\ܳ%[���-��DN彋閺~Q�S���%0'�b���p�$< �CW��\ �*G�B��j5��4,�5ZQHu^��D�'Q��;�#|���Ȧ�E
��g��Lc���."ZjeʡI|�����,\b��@����֞�6N�t\��2�)�9_�7=����l�P���Ѝ~��nL�bUO'ľ��)��r*:�BS���Q͓�_T5/��U�iE��E٢#(�������3ܴ�@>��a���n��T��-�4��!z�Fq��g�*���^C����cI4$������Se �5̸�[[X��o�((�q<���O��)�.�N��?�&�}�F^�}i������R�R���y��/3����/!�{[�' <���������W���߷ka���rs�Yve�֬xFIX�ش��n�.w.ޏ��x|52m�Hw'
�\ϓ���;sy?H��_���dI��L�p�K�yB��-K�d�?�����.u~�W"+�ڥ����l:g)<5��/��Z2TIZ#�z�$xό�#ƶ�S��o�����E�]( jK��{�n��y��3-�þ��dqB���8�,�p�(������5�� ��a��0)N�i�EXb9R�=��]�q��(lV�~��QO�[Z��*'��V�@�E�s��F���<��^k��A-u��� ��N��qk�7�P�/&)У�L�-��5�� 1A��W<T�� �䂓Qw��2a�x���p��tN@��Q��g�z�[,�ܛ�F�Y�������AMt_��0���ø���8��A��N�?.���	����qS漃^m$)2�7H0	h���w��S�ȢB�B���	y�2�7�m?�3��$��|b�[�_�8Ƭ�ŗ�]E�>����J*��<p�m�Uf�����G�/TX�����B��qP&	A,��N7��]`�%����$�S��w"1}%�[���z[ �>xi#�
����i�Һ������a�3f��mD���]tOh���ʸ-H*��#�]�0p�,m�\G8k}�kΰ+�K�o�5|y�P�f#�<�@�j�O�b@p 8 �5K��ѳ�W�؞�I�u*����Z��oE�X�z�����⎚C⮢�*?d1�i�o�ݾ"B�+��pE`#�Y���Ԁ7co�j~tWBz֌�
�����*G8��E5���q1�ߔ�M�ie�Ļ�2k��(�*�g�A!�x����WL�^#�I��M,�E@�7x����7.��g���)�=1���jͭ$cs�P5�n�]㳃jE�"�d�}����׮����guǲBy���e��s�#�bԟ��"_�'��=_�b:ͤi%+P� A��`��y�f�̮t���hlV<�>��S�ix$$�[ڴ��~��9�&k�l<�]�d�UJ��'̍�i�J)U��8z4T��i7B���c�ɓ��Lg����Wo}�qJGD�\�v�B��Cc�@�����Hg��õyL�t����$�$��M{��M�$�G���F5s�!�8�?��ɸ��4@� P	�B2�ߖ�p27�Q��U6�x����G���/;9��
%�Pc�� s�_��yl=�R���f1ql�VɶOw�c���Q�ؘ󦐎�D?WWֻkz�RqP5�<C�������`ې�J�;9�+�׆�]����w���$A�w�Z2� �<���]�f��I�bT��,c�ׂW�d;�o\k����v�4�V��K�����y����yo�P�����V�џB5N���Ud�ہɰ<�([��(Mػ �/���ӹ��z���*� ���j�eAi¦�9r����g:b��t�2���w{������gx�<-}�E�#������Ճ�߱+����?S}�+�T��ʪ1P�ЇH�A'�'���w�(��9u�ι�����]A����Y����	����.�	8���ՂJJ�m��-�x���*bܚ��&�ݴ��
�y����� �|&������D�Z��D"E�EU�Q-#ٰ���h�|Z����HQ��,�n��ҕ"8:���˦M6�~O-�1ؖ��Z���`���t9HxJ�T��f8Q  o�A��Yh�ʨ̹aV�w�(�n3�c�.�:B�Y$����2(~�_�9���,	���/�4C�'���巻�ک_�<�n5Լ%[�ς��!k�"���1A>d��(�ի[%���k9���x_U�ۛn�j�O����*����۳�[�{����0��tGԴ�u���&�	�âQ���Z��y��o0��o.6�eښ�_q�#]?7WYp�D�)�G�?�ŋ�.��$��IO���<%$����|��2g���<0�r�%�o����9�cr^�}}�YQa`�����y�x70������~�:��Mntm���l�H�Gm<��q�O�=��A>&1�7�c�@�[�����,�L1I���>w�D8�
�>M���*M��,b��0�ʠaJ�2y=]�x=0r��.�+�?\�2�-0ˬ;+���J�N�:!�P�i^]t1M�2�q�����F;���{6 ��@�8>����<��)�{4�Um���닟bN����vڎ�M,G����P����q<EJWs�i���?6�7�#��W��c�j���<�V���	f�������`LF@��<���o*���"�wK�K�G�&v��I2�_�/����͊��@(fu%��\��5&��7����X�Aq�2�C��#��1�&�3�
�m���a���&�`ۤ�Z�0:����	?'�ro~2���v}V'Ŝ��؞d��/��7�����p���� �ICFt��~��YRX�J~�a����\�I PN/��L�;��gE,Ԁ�͏���G��4Q�-��K�%�������dX*����P���J�Y�Rbώ��y�c�����.ĿH��䂉=�&�e����1�zoև&j�@���/�<�~r+9�����W	��P��\��l�pڽ�Z�~GԔ�R�p l��3xy���w��:�h����P�?v��Y�;ؘ����Z�4M
����PDҥl��=��_�Tw�MIMM�_��|q���p=E{;ܞK�r�Em;�_h4��'t;z�����)l�s���D꧌�y��2���%f����*����]�[^�>��95�v`x��h�7;U@[};F2�tѸ���m�\�&!s�d�L:h<ֱ�w	P`q��
��IJ�5�<�i�b;�>�ױ���<�o�:q6F.�S�8�픙4~{��7xtc��-��o�R���F�ߦ#t,�P~��8Nk2���7x*4������Z���֓�~<68��ԆT��׋�����оͽ�_ݫ�u���l��[��71���#Z<����0Kⱑ$
̢K�b�I��ڮO*���)�/�}�Sɧ�	��^KМ2�.�8���:�j=BYz/ qG�Q�0�&������T��d��4�<����%��"z���>��~��kB����XLO�Gڈ_q=�V/���'�X����k�f�"=�k<g��>p�n��ճ�+̝�t�-h~��3ח}��r�l�ay�˵�1/X�yo|r�m�F���G"��6O�	�5/��ZV��}+_+�`:��{?7K�5�A&�Q~K3�kH��Y3�8�X��)6��aT�r�ş_�nK��]���gZܩ=q��CQ�{}�G���*�>��g�ŋYp#~%�E��{��b�%@5����_�v�YЯ2�"U �t�q�xz����$陛�Z��]�\�<�g���'̬��v��ѵ^����y9}�V?�d����.�n7��|Ќ����|m�(\����j���8�A+~證��	�=Í�l�Dt��h�>�P��p�/�[�o�ȑ��N9[�HY�nX�x:Cd�'2.�V��׮�x����y�$X@拞��i�5�W�Z�%�/[t]���*�ML����R�&HL��o�5�j�c[uo����M��Be��~�q�)��&�o6���{��*���I���؀�H�R&�(�f�����K��E���s�]ʲFy�����AK`U��ῤ � ܚ���tX�n#<jw�aߣ��cn�X�o8�Ġ�E�[;΢_ř�EX�b�P�Q�$��m�~�����.14��c,�Y�Fr7�-auu��x�tZ��B���R�{�D��s#ԧ+�\S���NHÿ���X�8&U�;�J����\��Yƅ�S���gߍ�mt�����3�JaE�x�|��^�9.���\7����ht~���^ a:\�-q�U+m��D�*��Z[Ș��k����T�]�bTe n2��+�P?�w�b��8��&��N�/����T�Ր��[���FM2*�.�f�+uR�����a�*I�pc�ֽMF��o��J��H������KL���K@ط�F��x<�j�"_��*��L8]B��̡��,)�Ή��} ����G{�[�˰^`����k"HX�y;,cp����gf���[��\in�A'Z�~�+�������o����#c�Lٝj�s�C���(�-�7n
{�-�d�IR{�mǋ��_�y�R�S\io��.�Rt,)�;W���}o;�}h�!=њx���uՠWL� Iz�c��jS��9�ܶ�v���KZ!?�Kɰ�������P�d��u^IM;:?��z��<~�3�u��0p�����Pd� �o���C[;�J����<�LKP�A��p (D��?
��0��q���Y�K!�g�n�#ImO�q�/fێ�������]T�˸�`���jM��Tl
	w5�)�TK�_?�mͅQ �����M��[G��p�NF�dN���UtqZʣ�1k�n��/��[���y����ٓ�65�\S�DXßй̄]���q��d��-��	����+P�>�=X�S&���c��z�Ȓ�F�����I��P�oD�o�0.�X.!�t�i&Z�Bؗ�^���1��ie<09���w��Ϳwy�?U<��ۻ���x�6!���%�U�T�a	w͂����nw�Nh1�;��'�<P��I�|	g���j���ŏ��փ�YVڪ]�,���vL�FV�^�9��V��������w=\�y?�HJ_�����l#>�&	��\"8� �`ͤ��<(�D�3�li<�?u2{����U��N���Z��n,��R_9�6���D;�󯢖8�F'��mo[�n�ř VA���W�ʳz}{����8�K�D �0�������5��-��
ls��������`j�U�W{����βn ǽ�J^(�|2]t�~5�ECNĘ�-�l��+bv��f�S���m�A+K�w8V���,�[R*�t�[c �A�̬:�6͎m	#U��K]��׈P��v/��3�O:��5�� bp_�����;ؗ�a[��zfd�հ�QؚR�)6ˣaS�gT[y���U�,+��c1����^G�oU�D?�fI���yƨ�4٪Z؃5�� ��F���,:�GUr�;�5�Z�֖��脉L������J��'��nc��ǽ��?��x<��=� ����󌂳���c#)�CT�/>-{E�[i���Ə՚3�M�ll����̊��X��:�ź��ʿ�R�rj |�Ү��H%�&-xة(�nHF3�+���B7R��� �t�����'d�1d��m�� v�6T��=ᨤ�ݍ��ԸMs-*��M�m�ɗ�`#O}f�:|~�5��~Gc@v�;�E�c��^����ɿ�`�U��ʕ�&t��Q�(�>���g]M �)�[���1y�/3;V��4�{!?&#��=Q�T��&�5���IE��{~��R��@/M�� H�'�ё��½���J�+�e'��Mw�sR	�+�ʘ0�ֳi��7�����U$�Q�&��3�{��b�g"rtv4��,W7i^��2�O��X��gb�������@�:zqc]�94��r�Sׂ��N�L�+4��8�$��)��H<~䝸��c�X{�T��Z�	 ��߄��V+�A��X&�[}[�J^-�o�>v��D?�?򺬢�b2�~fWԸ�a��Uӛ�����d�y\H�12߰�d��Hel$�P5W��f�~1��f{�iSI�r�r-�6�ha������pm����m��4����������� ^>W,(���jJL��roH��Q�}�9]C_2��K^�0_W�&uP��r�����L]���^�Twj�����m<�-�����Pd;�k� ٩5��0���	ƀ���v�p�@��P&_b�+���c@������"�[��t|� ��&�A��Z��E��{s��#Mn헯*�m��WM�۷��22������s���k��N��KPbG�������
����ʢ�p;��
�����
�foJL� �F����bn��J�7C�R$������k�Z�p/����`!����8�w���?*�2 �����@����n�!�n���F�KA�������A��Kj������_</|��>{��Z�����W�Y������Ͱ�j$Y#�����������s���
����E�ʞ�;��b~|
P���DCB�{�MRO=L�+HƬ�P#��2�9 F��vt �ޜY����\�'��]�w�H=�#�S��q��Ym%#���'�^|b����N��� �;�a�;���x�Ȥ��C��~�R�|[��j8R��]�����Ť��R��8ań�P�]G��Wl��x]:#4�̟5W:ē���M�rR����m>Aj.�%ME���U$���������Qq �d�s���j�p;���p8�����=z�uc;K�N�|^���W��pďJ��)��
�������=z����a��6�"���w�f�L��o!g�i��Ӓ��?�E��_�m���\,��8�2f�@j�3���I��@h�8���&ш��0|�n
9v�Qڬ���$[�-��xK]���/q|�Fڭ���n'<���B`��- ѳ��:m����Ӱm1)��\�O�k�<��,n\=�.�Þ���g!(_x��"3����]��=���&�oY� �5ۘD�	?1�'�#.�f>{;)%�ĳ)XH�ǲ�4dcg�׭��T>�5LH�o�j�뮲TOi97�n�3���7�O����ĺ��Y�h(A�(69j;.����5X���n�1zl>4m ���IT��\��/�^#��*�$���<}��'��G���nJq���oǍ`�:(d|3�Cu����?��CW��vF�Jˠ���Bw�#����c�����C�ϣ�z��~7pYʧA�0�A����.�^�Y�Z׷-o��G�T�@ �V`���g���=d�o�snb7�� ��� �ͧRe!�$f}�j�{W5����t�����y���T$�=� �e�(\V�;b	zMXA]�������ϿbO����V05g5�n��8�W���w��ߺ.�X��f�&�sgQ����s�������+z���,��{�ʇL�]�Th�D�窆Av�Od��M���<�'c1��X�t.N���Ѐ�f�X���Ry���ד�>G�KÉ��Zk�+�d)�"�bY��Q+��jYR~�t����>��{}��>8?��#Z�yF�GU���;���~�V�z���9'�"��o2�n}��B�������Zg�7s>tT��-�
C&�H�~6��0ϫ�`�W�Q_"̣�$h@"�/��ꆕ��)7����L4��g��[�C"�K�ϣ�(�|S&�����{���t���q��_���B��`�j:�Ȏ�x7�'"K�s�cNU���F>#�����y�,��*H��@�0a�	��k:�S9
�s��_^��]g��fT�yш�gE%�5n`G�g���d�~r5^]`�~��R�jEzV����*^�l*b
yU&��M���C�ۭfcE�]�7�$%g���e.�����Jp6�t�ڹ >�t�1���_�y؞٤�f�͐�V���Ϩ}]wݥ>WAZ�]��)������n�v��M[ܠ
בt����}}\� g:pk�$�{Ȧ��xtι��S0dU���ML�}]b�.[G���f���=��h�s�L��K�Q�^��q�]�����x���R����;��1�c*&Րǥ�������+ϰ���V)a+W!�z���jϰ����S-}��f��nZ���⍬��t��G:�Ò>Q��*�g���:��h�x��;Q=��j���D�p���[r%���e�F�q�ם?$��D���D߬�q�.�?3�΋�7^��ͳB��|�\�S)�V�%��BЧ�G�D�7��i$���b	<�k,�����*~��9q5b��'S˺,�����q2��k��_��5�1��;����X�?'8�i�$��.Ʌ�l�n=�ε[p1`��J��U��3_ىm����t��ԛ/����<_��k�o���4��|V!X����2��I>��ī?���ҍ�q�fKѪ�1��JG�Ʌ&�q2ϟjR�]�ۿd#\M) �5�	��t�2g�l�����G����eY=�䟌Cm�מl�0��sٹ�$(J�e�X��{N7��Ԓjӑ$����\6Ț;������^�kh�W�9���� q��Nq�]���91�k�a��w�����Z�ɬ^9��T�g[ź�D��^[]��F9S�f݅��v3����?j��|G̾Ux]�
R���9�6v��0yd��
�e�����2�J�Z�����였�܌�pSP-	�
&��yݓ��CPT✴��>�#���f3�$�~.�qh_ܬI�c���a��N��\�bo�z�ۛd�T�^E�o�1�\[�1��yǥ�����*�D0N�yG�~K��6e��(�t����m���;Nى�GJ��f�NL��W|�_,���Mϝ��é��p�R�ҋ;��X~e�ĕ���P�`����2�@�߼{D4ҦN{�����M��CP�
U' ?�uxD���s5��ĳ#�raq��5�s�~LQr9�`<�� I�{R�=��@<)A���%MO3p+�ۻ�y�'�(�`��x�[F�C���ϴQ���k¿w������m�����K����I��/�0��G�d�.�� Z��ݩT�	����h���K?N��}g<�ֵ��61]�b�ᇦ���p��y<�(sdY��kA�C0�����52c%g��DznЩ����d�Ә�m��Q
m/E�'� �m�pYB(�蔻{ᣇ�����Pp�n�����m�E�f�>��,��?�阖����\dhp!� ֻ�0Y��Z��r]@^���|�3I>�}��z���_������a
.m�>?j�<^v�~�*�y������ʋ���#��x�^����Œ���~���I���F	��|&E{O�!�������I�T�a֢�oK���O-�r9��g}��_�f�j��.���,eN�3���,�\eLsdvl�af���0�3\}Q��Gȗ����.{��[�x�HkF�U��br�~w�<`8�}Ɛ~����-3}�� 
�e��&AÊt�(������N���<hZ)I�=���pٝF�˞������	���S��������jdP\��1Ҹ����	W�U5n|L���������'b��l1t�x��Ē	^��3���<1tmxY�}��GDc���@���e/�%_�R��7N��)�3U�$x�Q��C��P��K��0��QKp|GY��i�w��A
���Ku���Jw�f�&��/�Ӹ�ԕ�S��U�X8��<����S��S��y����j��J���'��tbk�B6X�^L�1šY�)LVJ���R�����Y�����K��wdp:OF
�%�Ri�5׽����b	q	���4���Y�}�c�.��!^h��ܽ����z:fס�,˅�}�ثW��r��B�SB7`��c�����zǀ=���yy�5�]�f���K�n�}���A�h�*}[�L��WU>�{"�)�� �oJ���zk�۩s�̸���@c.���}�|�z�&ߊ}y���29���G��%k{� ���zJ�#K.Z��Ѓ�]<�Z�);���Mj/C5p*З���xs��y�Z� -���mG�]��m��l�8��nz���~�S��X;'�����T��-f)C�;\��Ό��y��{Q�W���� @�b�ģ�BK��*�-�1J�KҥV�
�5��_�� V2���5 �]Z��SJ$�~�5S�<���]cre�h��h�Y1K(F���3����i�3��L_�>�P�Mwi��#�μ�����(]?���`/4���T�\T=6k]a3�]�{Nߑv��0��ۓ̹��"����N2���!qj�ݵ��Bp,Aռ���rҫ��KR\�4*1"d�֜Xe�����⽸�ڳ;���e;����a:߳��������=Rt�Z��$:�u7�e1݀��^2Φƥ���I=XE����L'��Om%��5fH�k��K֥�fjtz_�y�[<�I�jC��",��0ڿv���j�-��./`�T �' ˺��9��S���N]�u��Fv�U�/�B�������
���e�g���	`��ɥ��=����+G0�Y����]�&��m|�d��8u��J(.�^�Ҁ��SDJ�e},�]Y�J;*k��i��`2����o7�B^��"���w-�sI��_��l���{K)"w�R��|(�	�L�/�lM�\��Y����6
O�Ӱ��C��,OG�%&��/��ؐD�bzZ:+�fH^+*X͒�P�,�����}�Z:�I��d �<�ɴ���/-�Y�/��b���ϼ¿�t�SoB3�$ռ�y�z�6,�9��<�%�)F��ߝ/N�u��B�n�S!ޤ����aK��ϐ|JI�ooMN���D�b=H+s^ \ض�e��,�sA�Ӯ��^��$�1��'ɑ�q����M$_��&��@�-��"&rw� ��Ʊ�\Er������u
��\ �'�����˭ߦ�,]n&��M�6�[(�,�r)\9�&Ԭ.�3�)b�`V}_�G`Ɵ��׵�D5��9�7��vST@Nkm���k-�T�[9(v�6s"���Y����׻��۷��=�4���$���\���σ'~2��K �3�����"~�� J���/��h͗Z�ZG|U.�e�������G�g�Q�n3�y�֥��#��V�ՇZ��/��_8O֚Y�tN�uq�+��=5��(��]��l9���L�|���u����r��U����3���
�~Og�L
��~�X��x��N}�i��@b*�6�s}���G5���(L�>w�|(�Y7?{ޤXw�!�ǿ��c��k���s��R5P�Q�`��r2���w-�c��!�ג�'��7i��蛘t��J��Fg��x�M�;�~�b�����ŴyPu�y�#��ۖ�C�q�NqM�6�O6�D��eX(�L�\�ж&3��Z|<7��3U��k�m5���d��V�+�*T���1�T��IM���@n�}Z��+�bL����5	SN� V Q5S,u-�ǳ���,��Q�_�"d ݹع���"��hy��x��[�=^�r��]�{����Z�P0%U�y��p��B~o����~�o�#��q >%�u��<��Xe;�tc|<�4���=�~�S������)�9�s�zC��I�B/�(�E��w�f�[0���3`������8����䯺��5.����9�N+�� �����P�=YN���i���P&��?����@�I��r����V�`���&5k{nӱn���r�c4ςfa��T�!����,K}	*���&���c�נY�&-����a��=K��<G/����jӛ휈g8��@/Y�N9(6�D�Ա�k��>!D� /C�QѼ6,�ߟ3nn�L��3 e���n��spk��i�>g���*tYl4�!�$SͶ^���y�e/��	�����cLFk0�^�BvI�c��>�㊽H
��>w@'j�1�埻��٪g����
��7�����Δ��<���O~j�������%>ѿ(��V��Y�m���#�#�,��ؒ�~|g���Y:b� Ǩ����6g";Xd������v���|��N���,ZQ���U�<�v��v&�Dϱ\���z�x�J�K*���"�W"%�K�x�^:K�pv��b��mݏk��T.��R6���Z氪BAB#��²���\�}��9uD�Q��F��Z�G\�_�
E>B-2�#�sO(�=�y�	�}.^�X�p�^��Q�y,�t��جT@��X�\z��[��A�샌X� j��4!���ՄYM�4M���%.��ي��)au��z ���䈠�~��@����d0�)G��d3h��H���{�M)(���4�����Z�E�/�,$��xG�.3����4>3�GF�0�]� p,�NVn�	�����CA��[>ޚ~��N�w��G�*���edt��C��vk���a�S-��A�;Չ�z��~NMX�1]��D" a�r�d���c���O&N�y��<
�y�R�#��l`z&���-a?݈����mH_��h�Xj�M�%W�Y��h}� ��E�ofP��bx�"��q?]Qc}��<M{' x���_����>4�$�7�L�?��	.��z��	�������q�W�D��\�H�˼��� 0
������cA��п��0
@45�H���R?Ã��b���Fwlprr$F_�;L��/�F�/8A��j������@�#$��\���o~<X@ױK�2��� �m��*�q�e��u� ��8�Xը��y�n��ս�2��:d�B%I�w�p����o ����au��c��Q��.A�7����	S��L'x-eq�[�u-�y*��haV }�U΁1�(d��>J��~ӥL���������_��U�)G���&��5&�ʹ���.��$";������B�"cM��}@6g����R�o�S^ ��H$�x�<~�i���#ӥ��y����?�W��z��E	�S]��[*b��$د��ҺV�k~�ˌGQ��S�J�B��PA�?2������al�l��zj���
ּ�<e_�?�*��*DZ�k��%aI�ܘL���'i�t���SԤ���-�l�#݁[�<cc^;Uf�r��!~M�|N�����X���{�cZ�o��-�c�7$��-6S�e`��%{��zQO>�v���%NX�q)�x�`v��@dSc�_���j�Q+�m�G]Rvi�L��PZ�B�=�YV����)���c	{n8)�Ķ�C3��q�?�F�#�﯇�*VۜXlzf�	��:,�)���T�?�h�eD��%���}�_�2ٰbE.]��2������?h�L���l\�v}��~J(��l���\�ϑƩTlP>�$\rhı]63��y|�6�"�@=v쾛�#���"��Zk��:Z��#��H[^�Ӡc�Ep�AP����_�z����l��p�����i���.Ky�3�?,|�"�b����)L�c��.Wc�����oQ��2ƽ�7*2��;�1V>�����;9��L�@[���&��ߛ�/��_}1�ϝ�~����Y�����؋���ķ8H�
���aDΫ�v���ŵ(���9x�-��l������]�>lG�ZN�5!u�0@�ٍ�Wo��W9�=��A�5�'|@`��B�[��p�7 ^��d�&�y ��R?#�|8l���+l��Lj��2�vp��fkyλ��
H-����[�_O�22��%l?
��@4b��������W��ҫ���-C��'}���P�mKZ��]�0�eX+2���SW���e힠ď�P���y5��,a Ф��g�o�E�X���.:t>X�c�<2@N=�*%-�o�RL����#[�E!IW�t�|rH l^
�4���8�p�:^�e6L��ݶg �@Tz���\<IE�$Ie������ؕAD���yoݛ?2W�	c���n
�5�2�8�r�e>�f�����e΂%����]��c��[��(qx��F�fr�����PǴ\2ֶ��A��� ۜcg��;�������*���h�� �@R�J7?�X�og���9A�^Z+��M4�դ�fQ �M7:]�M�/H�;U���+���c�]��7��\mau�j��h`�Z��D��1���݋e�q-��RL��n�1LY�%���@��C�P��������@c��s6B�ש;�e�o\��qTW�vߏ�V�x�X�CO�y��F�]�O^(��ܯ%h��bi�����Q-�n��P{�l�*�"[���v��8ӧ6h}��\'[�F����ާf"r�=�p�Gm�41�n��H�W?ſ���F����[	oy3�w~��JI�Ϡھ��(��{�K�z%����^�zU�h���� ��я��Z�Z�+�16\_�9��Ž��&=A���xSw����������t��>!N�T|Z{c�~�ηk1p��Y^���$��3<��q�����9����M�ѫ�������\�-7�h��;�e���ܭ�A+y�&W|�ۙt�������K]B��>-���ރT�����z�l���E�Ie���c�65�m͂�?��qx�E[4��{�P=V�5�=*_���x^@jȉ$��z)��"'�='u�/��� �6�X�q�����Ki�>�����pb}���GH����[)P�м��#�� �7_��@<;N�sh�䳩���ǃ��g;�[V�c�H�bo�-:�R*�K'y����w6C;JT�Qv2������}n y����1�3{[��S���P�`�8K��E�����s%��^1Q�E�����f�Wci{�b��فvE�z�)΃���'Fj�,!�EjϨ�#��M���en��9#
Čg?=��um�%��+)�+ۡ�Y`28@�ro�� g�5y}^�?�Jq2�:Ʒ�߬�%_$��Ȗ��-B�"?ÔP\T��!�V�I���8�{��xn���ru����>C��ng�i�����Z��;[��>�)B7 &�[��A�J̕�y>�-�E��\�������9&!�f��|�j&ڽ�_t{g���z�3`L(�3�um�q���@9�U�Hqb�z�)�d!;Auo��]n[�&�IR��o�!?L�(�����t���jM��i7�B�#4���r=#�w�kan�q�@�Sѣ����F�;-��v�����q�K��nf�����t������k�N��d_sa-�25=����?�'ڀ���I��#(�La��<A����_�ξl~�츊�z|7t�����y�#)l���:���[�{�^3յ�J�]z�n�
/[OU[��+����k���J��_�fh�1=�E��(Z��� `W�V�M��Q��nrj���s�V9����tPy��p�0��&F��m{�~%��[M;�iJ���}�|d@$���r�V<p�����4�f٭���	��z�jm�o�L���t̝����|O󱲐�{��TU�����k���Z�-�J�j��0�f�ctG� ��z����T�I����z��>����K@�AͲ���	Z�y�ͭ���hIkcO�@�Tsl��F<?XR���Jw,P�tSf�6�x�NƜ���6n�cYQ�A|�#l��~���4������ �[�e'�������:J8=2�GRJ��e�w�;-ݜ(8�웰'���@ab�̹{���`�#���5V�לw�H����/#ʖ�[�����ֶ2�9сS��&��"�����:�ͺ!����8��Ҽ�.�WZ�"G�9�ȋc��bƊ�8�o�|���\�牢�� G.(A�ȷ:���li���WA�W�Q�R��Q�Kk�y��5�횑/��X���4����u��[_А�����}螥��R(��?�r��e���Xڏ�����,�I�Xשt�]��ϗ쐖�F�~�	RU����b�u�����<k�W<xF� 2H�]����y���cg�6�:$D;B��q��(�p)!_�X�&OMz��G�4���ͪ�QZb2c3$g^8����>��q�G��fQ���b�4����ziE����f��5�&��,�I�h�6����_,|�y���L�^�M�@7`��艹?䃱�J�p1�?�����)~�8�:�~��2D}���>)W���Kw��s��&��
�iG�;K+��E�OᲒ�[���J{|X�oO2S�7��w���#<۶��9����dpL4Rf��5��(,���ۿ�����GwGi��H���)�uU��D�S��x,�����T�6O�s�����\��+�@%zF�3�{�(��w!�	ݨy:�+�����H|��\�bX�v�7�`/C2x��9��V{��%/�3m�3��i菖{��݆�&2Ci�!�#��d��{���'kTu2���[r���@�x%�G���	l�|n�ۮ�p�>��@^+�b�\�7H竎
��-�|M6Җ��z��'���- R����´��i����ﻗ��f��#�$2��@`�7��?����}[|2�o�p�^�]Y�%T�Z�7��[��o��3�O�'���o��K�j��"iK
~HJ��?5N/Pޤ���MEz���৿O�� L��6���$�ǃK�jR߽*0�k��P/���z��e��CM��G;�WH\>ɤ>��;���,Ǻ�^��_<�&_ǔ�'�,[!}��gI��,i�I`GД�!�'�pE��Z�p.�3���ٙG2)�F$�3v�6����5�}�*
l��4_�c�5/h qs%��MPy}y�Mk��^���IӤEv�m��"	%�P[�9n�W�F7����A����*��I9{{:W*U�o%!��ʎZ�{1>HCs*S��|�fj��Hzo�(p6�9eX���6B�ܨ�X�Rʵ�~X!y��f��ާ��oD"��2+J,ↄ��Cя-�5[X�3�y���D��u����q����~�f!ۓ%سc�|mm���֞���#b(�]������"hlE^�|��D���{��Z�x�!D%<�9��i�lӳJ龐������W�ɵ�7+|����
M�,�A��iś	�����E�f{`��k��T1r�ʨS��ȣ8�xRTIIɺ" ���rU�����2`�6_� 
�B�<�Dd�9I�`U%��Þ�L?7Tk�On�P0/$K/Y�����#�~N�Z��K�v�c���m����M�(�ʀU��,T�˷�ly7���)���[��� ��)8U㴇����t�^�X�&�j�\-��a(1>�F޿�}��M{Vi�U��G�	'~֒5�J0@bo�s=hi�IU�I)������a�/��J��7��i��(�Ȁ����)��]$�]�wѤX�{��o�L�0N���+�^�܂N��e���T�8�����n�XQX2��j%<C��4Э��[���2e[L��L'l4G-r, �le�D��0n�$�fI7cA���}0ߦ���N�#�s	����.@0�rg �0���R����V�ĩ���<G�4�qG��ޘzj\��.ɡ�Pp����>����s*X���I��#]h_������G_��=��3�$�����<��+5YH���)�t�][o�4Fz���{v�uIs�G!{y)ᢱflŊKJ�����+:7� ��	'���U� �+k!�Ch~Q�ҏ�M���V���a�O=�أ8��alջ	�)S51ՌÍ\�է�h���H�x�+�x{ =��K%�z]���l���Jq��>�B
�����nz�m0R7HD
L[?�\�w�˳.����SחGz�~�%r<]���>e������L88����9O�C9�(W��r�RO�$�t�����U�ͤ8|7'H}��! A_�8��#CǨA���qӨЁrO`~F�es�&�?���J7!c�Ⱦ/�0N/�7��s,���
;�\�#,���jeQ�������znxT.,�K��W�R$��
�6�"�)ppx��Zv�*���C��o�Q(��H��į��6�x�	0N�'|��g�;�!�"��d0��N�2�'9J.��kl1@!����c�ނK�F �C�9��GV��D/+`q�
��)Y�o�W��[*M�}�v�*g�3{;7������@!���DN��H�]LsTe�_ݒ���'����L�����d� �e���DǮ�0���2���q\�ݢ���;�����3V��vo�@��$��b[�K0<���^x��-@�t_֋[�$o�}�㤊ݕ��k��wרR ��±�D!_&R�*H��2
�LQ�n"L����D�K6��D('��?�\�[H�9���^�bL'y�*yt=F��}j=?$������yRnMЕ Q�!������5{b�Tآ�r��Q7Y��>K�ݪ"N��C��?�#�^0��Y�HKab\ud"�X��\�)��,^���^0��	�q*��d�0�4|�/�CG��޺���s�N�;�Q� �/BL?�!K`6҂��E��]�_����9�?��v;��Ȍ�2��0K7�d?a+��`M���,�3�q��~z}�'@������%��k��#�^oE��5k2��t�y������mB��f�IIw�9:n�|�2�r�Qh��L��8�	=�={�(<�؏�ȜVZj� ���moe�ɷ�+��s�Q������	��>��R��4�=2�1*�|�.�����|b�3�ף�D<[qO(8�[�Q��j��ͣ�O�U�{5ocv�H��Fg���'�	��� ]ҳXE� �ȷ����|�(��!����F�����
�c7���� &k&Ι-�<�%�M����l"��Y�7x/0�"�>�\?�*�qE+�1�![�ϳ��l�AD�R�5h���n�L5(1޺,�6�<17��W�W0YD9O�i�1;T��0
��Z�d���:��\ܧ]~�����b���S���45)@p��>+� <6@����r��r�28��YG�hɠ��9C�ecCN���"�3E|_y��÷�l��gF{�}�=Lqc�H�o#R�cF�:���{ty�������b�����?k4�b��*�諳'��t���b�q_�y>B�Qx��k�bS�ؒ�]�Z/'͜u�oJ��V�i�=�T����CaCav�����G��֣���l�B|e��Ȏ�=���'aF��>F���1�/��I�o�pI��N�J4/�O�1ј/���ᑔ�]?�3�b^��Sip$��I���Kf�{��>�����\7���_W�m%�e'$8y�����}��~@īP��t������^�^�l��o-���W��և�F�Ζ_�����z:s�^�}�#߷Xc�<���T��M���:�J���ڛ�ͫ��/��w@{�������՞!�h��**��x����;��i�����n>�$��v�vv�P�!�e�����T%�&�����k�N���;ǒ��g��o$���1"��'YZ���5��|��]����T��%�Cl�[��/�������32u�I�C�qM�V!׻.<2�˵����o����C��|� ��e��|KJ�%b!ݍI�����r�3���������慳:Ֆ���C��	�2=�y�������A�P��g�����W�l��p��1|���Ȍ��s,����Q�=�������ZF��f�8�:���KZR����QTX������֤Y�r�]�TՖ@�����f���o:?6�QiM�$�e�y��_e*k(��ǒ�(υU@d�K���7L߲M'<.�/J@��Ϋ7}������\�Mh�@�j��f��!쟕�( s{���RX�*��ff�ٯ��P[�X�$��^�Оmd<�^q\���d�ɟ�m�5����T#��F����ظ
��O1��� ��ɓQ�x���L��/��8���,�0"1�n�z��jWXVf ���9�hȜz)�GYqw�����ƞt��+��� �c�ƲSŊҬ���A*ϧ�k{E��0+�5���$���:�D�Y�,��g�f̲֯��w�|U��'�m~�Œ+1���T1[��z�Y�kٸ�=��Z���UN�s|UѽVj&���4Z�%e�ȗ3���.)y.���rЊ�>�j�nOR��=?��/���BT��p�>W�?�Y�v���^EķU��.諸� �܊�g	�7�~JcG`P�ʸ��>�Ё��k��ȧ����.�4�k�<"��; [:�r���s���0��@�η��Û58��4W�B�h �#%�K"�4��+՛��BV4���g�'༈��zs�eHu+�/!F׆9X��� �J���WN�+@����y�taHtI�r.� x?�X�(A���vo8xG6�"���P��@��/��\�;ټˏ�},U,)^\��_wL�j��b�:��q�fL����]����S�xμ2s��_c�	g�k�t�	��
*�H�9�#䑏��IH+Ƌ�����"��>�y���aK����R ��xD�zG�BKF�q2�@Ӌ�.?�'v�I!��@�P��6�b���6'+_���qw�V�%��h�oR��	`4`�s l�|���L�m/'ӿ{���vٓ�TG}��`����&�x>C��t@��g���z��c��� [G �[R�|9<��g�Cx�/�y��U��잰�[r�Is��j, i��zіZ�Q�8��>��'�*���O�%q�k�n��J��BY!N�oC8�I�gut�Y��!à7`O��p��M�g|�\2�3(޴������P�a8��t��8��w����;���3]��h][���N�Z陘��	~⻺9D�M�	��f��I�������@�U:s)K$Ÿ��z9��7C��8��6M*�T�ł)���Kc�u��7�@m�wS�J�6�
%������/�!ׂ�=Ck	K�ޥi�9��qr1rϿ��]&?���;�����ʭn���Ao��jz
�������%���k��9��˷r4AH^�;�lO�@��8O��͢����$@ҌvC�QhJa�U<��찈��~�eN�{�E;C*�:�7�ҁ��(x2=�����K�KO@_&$j��z���5h����%�����U�v4� �#z���h����ѷ�s�H^ThB�wh�&���V.>(�#Ӻ'�D�[qVO$�Zk��'9���?�{@
E;e<_�����ʣ���&���G�@N:w�Н���j�Wd@foNW6L���~����J�s����\�զ�V����=ʿc`��#Xy4�f��!`t<s�끏?"S��Fy����ݒ�lJ���_TEJ�I����0)�.pc���2Ȧ{�N5e=/�d=�� ��� D5�1>Vw�s�����;E=���IF����3�W2��D�$k֟��:������U!+.@��s�휰���V�Q�{�7,J9o <|�Z�U���:o�Yy.� 헏�н��d�~PBt�tt�rt��	=�{��c��<��Pn<,U�T�}W����:����@�2�q��w��5�	|��2w�=��E���.$p�Q@�
�UUx��Z9��x>'�{�Z����D1IbJ��q�Kcn�شj��QT灜�G93��)�� �迸K� �2�v�;�$��[�xpL���|bW�o�{/V_A��Z_���C,_d �����K�}����!��q�)?�b�C�y��	�� ����ԍ���n];9&��n��4�N�(C�7��n�p��hK޶����r����h�������e�zڼ���5qb�24���Vh�xM������(3���e� �!/�&+�� � <h�B
W=e�:r��I���iD�򲓟��a���T\_u
$-�F�)q<Sh3#f�<j�Eȹ��M �v[���#��f)���\����Av�}����D5*0��3�0�%�L�����Q��FB�'%��dqL������>j��:�O�� �2�X�N2YS~��*��+�����F �[�ͩwx�MT�p
�	w@��QI<8����|�Մ�Pd���֭���� `�(���ՆA^��.N�6Q�rs�������xm	��)�Rmc~�W����|���[�SeA0Ё?�ֵ(��A�d�>��Qk*��i��EL�eb�@������_��]��U�Xo;x�@��W���Z}��jT�E?���XcA�4'?-� �yΛqΞ�=\Ē�
ݍK�r��0K��l��p=��}�D��M���5F�q�9�ر9?�W��'>!/����{��%�F�0�3�*��Ŗ������ܜX���dJ���8�(3`�z�d�MznFA�H��� a��,6��U�>�K�]�l+��q�Gl�n���V�D5D�+7�U�%��;�?�Wp~�����ZtF nm��ye �)�$�\��b]�-��1;y���>�4��t��������5�����Y�
F��z��g�m�TH�E�q�O&���~��"�d៰dċmy,�����F����X��5�����6N�p7ZO���9�.�革�L	�gQ�bzR�&�^X�O�G�up���/��T$-�N�+�9^e��|��zs���K{��x�t3ﲐ��O�Ӣ𤼍�\���5�]K<>^��
�˓Ά���CZ�s�� "�?��x�ꆎ���`�m]eW,W��F/b�=�#��f�&M�-��~_��T}NkPCJ�C1�#l��kq����Vc�K�v�0�\]8�$]cJ�J�Ct/hq�l��0n�f�췤�VɼI��g�,��A�1z!�W�c�;b��a�F��>���ɶ����L�uK�3�Ft�e�aTc���oV&�SyY��8��_1Fq{ې���xm�������D����u3��lI���%BD�o (�~W���(��+��2����SW3��q�>K:�� �'/j�v~\	Z�O���T�Ѿ���������y��� ��SǷ�T/�j��җ�(�N���v�U-�n���(I�ҧŎ����x�]z�W��|#��F��w�4/� D]߽�2�s�!*�}�_�2�J����2���E�#<.D���|]�D�\��dN����
�h� N��]&�&4�O����Z��T 8�c3n������l�����u $rxj��Sv�m��!���C�J|���3������]n��ƩC���%J?čO���W��=([[��p"v�C=����Ϳ�۟�ڳ��3���Mý������\�C�ǀ�J�7�+�kA�iLi{�lN��K^����Ѧ"�'�C�9��Qƛ�����M��9���B+�`x�75��7ļ�#�J}��׫��UK7ͬy7:��?��;��5����E�.ME)ҥ*u+E�
"��Iu���"5(��k@"]:H�P�$!����.�������7sf�wNf��k������=�"��o��M�EBMT�[�4���h�`m�e^� }�yh,��3Lu��g�}?S����]>����,a�O	|1���j��Z�����"Y���3�?;Ǔd���gh��1���k*�:��d���8�D�����tm�Ǭ��h����Ѧe��t��*���'W�<�J�j1)�Y!Q�)�,�����H���ϟ3z�^sE?MPnziN�(P��J�}_-�'� ���jc�(�/�p~��_�\���?a�A!�;H�|Zm�2���|�:�M��<"��ۦ��m��V��+�Q��S��w��~�a_r����w�M��0h����9�(���Ǆʻ|�Պ��O0[�����vM��>��?_4{T��i�٦��8�[�>c{��tI����=��E��ڥ�wP��#?Z�M����Vqj��i��ae	���x�"�����
H{8i���M%�Y��)wǖV��_K�'�9H�W$@/n}`���=tZ}���}���
��[��nO���w���jşX�
����*��K���+J���>��2�9˽l:��qv�~�Fk���i�]W	�x&a����Lu^��#����%��++�m��y:����,;@����4i	&�&w
�},D~���>��[S������OAZ��x�-_ؿ�6?fQ��i<����!�L�N<PDȡ����(1˅�F%�zO���Zs�n�W��}��J-��؈=°����+�<��mD����`��0n#� ʂ(W^���F#tLh�é�Ε�13��X,�m]��+��?n؁�U�'Q
����p��c`tijG�-3M�|1��	�:��:!����䡁<u#O;���H!�
Ƴ��u/;�U ���h΁E�(�0{��g�]?W�>���h������/�x��iƒr��p�z@�rP#�_|K�D���_h���E.}w����YK�ϧ��7 A:�~�2���,bⲢ����)oFFޤ�n�6Ƥ�j�W~�g�;3��G���U��F��h>��3I��H��vn��Ʃ~�O�{h3O��e��7�{�pW�F����'��洈��Ÿ�?��3#�^��w�c]���ɯ�s6�܍��6?�:
;�h���b�Q�"��f�����a��x����L�ia�������)��L���������=ZO�i.�^,�7y��ڣGS�f��G�%�]����#,U�j���ɎQ��0��?z�ʓK�O�t���7i��T�'Sw���p�?xS�:�R%=��'`��?s���E�Ȗ���%>����d#o�{�7�=�H�~;b�ݧ�
ٝV��n[4�@�h��(V��5����ӽ����W����s*X5F��Ge�Xܶ���N5����`��|`)�����6���lxֻ/r<30��Y�-2βAZ��o �&E��?���^�_�m��>�\z:�j���DY��	�x"�s^��4zh�m;%kz)n\����Ҹ�ҧ�Dݺ�ú�*��m��<v���P�T4و����&�q�$�����~�����4�sK��P8/^R�}�E�������ꥴ+�|VӅ܏S�I���Jy;p@�%��c]��`��'�0�I���m��h�^�d��:��v��vz��ޚ�[�|6t���o��(�&o��KKm�#~=�>���^>k_���>:���%�:_� xuG�35[S�@������&U�=J�G���pM��{B�i���W�՞LyQY��;��Bζ�T.����7._�֗�en]����d�͟
X�J�]建���E�}�����2q��n�Ӓ��w@�t��D���v/�n��=HnI)�d8X%��#�x�>�W�^Vu�w�ӟW��P@����cz�"��|m���ő>��Kr2j��@	��s�x�Z3^��w��(Ґӄ��<����ːr���,��֍�˕���l��V�)�E��l�-%i�d����q�Χ��S˟�����,9�����!�8dZ��GxR$��e&^�u���n�:~�z���J��H���Z�NB��ނ_���lqly���6~kE:�y����з]u��8�Bί�h��p�1	V��o�/i���y�D�Szc#�����+���b��;�(�N�����~�?�ҭs�H�g`�����&����b7�|�X�7ϴ�Zb��PAѱIA�J;�ZC��c�Q�z��w �qޣ踉��Xʍ~�G;F��K�X�wE�<ӯ �0�a�� ����@�#���?�a{�֞��ŮM�yy�c��b��^���|���qm+�a������ƣ����,#������S��d�b	]z��2.������VR�T��͂��E����8�J阗� A�r�q�H�]R�->R�$���w�["%⏫�'��k��ҧ��Z/��YR�ղ���θ�.	|�W6`�.ߥ�����;��}��"#��fG�g��%	�:b��I��7Z�j���������r&�E���o��	������O1�b�&D@�J��p
��]�E>��l�y5HtW��L9�^r�͖�4���>��^%a�=�f�"���?�8
�b m��Μ�Q��J������͵{�;�[T:�M�5/�s�r�c��1kl0�N�Ly��Ґ<k)�N�d�~h��Ҽ9�F�/{ta-ݼ?�k��e#�D���}}F�$��\�o����|�n��嬮|E�αQ��Y[s#[[�n1�M�}7�=w�[ɱr�y��C>#g�RC�"S}+���8�&1��������и�F7�8/W�,�`Êi9��6�A?Z�7�Fi�Nx(�>L� ��u{HY��(��toJ:�=6�%P�<��4�TF��!'��+�??�`�A��h���ȯ�ɽ�<������p\M�^�；H0 㙟H�zI��A	�N�^�ia��R�=��'k�8=\Э�ߙ(y]����0�,�~)�O�גH��nC��ZkRS�Yٍ���D�i-�*��ٵk��M��4�����6�d�:�~�̂�!чS�yڲ�˨���T�i�={$�+?���g��㷄���[��m� oi���>�%�4�$9�����N��r��6���\`����OF%�k���g�b�~](��?����
%-�d���p�I>����_\�Q��x}�����pTK��kI�N��y|���@�$�g�_:u� h��O�sY�@>�"��ո��b��3��P�~崨��ʋ|_���1E�>��k��}	k�S�"QUtN�I��_?{}�). �@�8,��ۋz��Zf��yd��k�b�䜧�sɩ$Bx�A���?zHq~?�Ҁ�����m�b�I��:�~q	�� v h��b	�US�����[1j���(��.�7�G~���m��m`�P�d�V*)���/mT8o�o�j'�e� a��2�G��kE��q�1���(!�Q����U ��g�F�;c���.�3/7�w���K�',��W�WK�!;wg��D����h��joCʇ��ɬ���>Y5R��,J�P�G]�t}��=�{�8��P�#n�JY�J�y�~�C�СC�I6c��zS�[�zۡ�Q�lX�k��!�&O�b�k#�&�w���6�V��
�iݲ�~��& r���׍2�5�����g%�.F{K5<Q2�w�{�{)��(�2���el<�H��[}�F�1�)���Ek7m���&�$=��hY�}Ky!,eU���U ٗ^qv�	�5�bk
v#�	Lt��Au{��icF@�ۭ�h/hnPD���M(����&����	��Tvnx�m2�b~㜭	n��q<c꘤1W�n!���d�Q��y��"'��Ը}�μ�.�ZB)�0⋳��_ġG˻Z5߰ `��(��5����h&|{�r�N��i��A�L<��P�m�D��Ź�ut�"ʾh!��0M��綯9���E�}��i�FD�ٓ�"��E]k�J�p�n\q�3e�GL��ɦ��m��o*{g�ׄ�LBi�.�[���~]��cޕ���"ʦ��ۦ�SL+of5r�<҄h��k[v���:_ؗ\���4Ƭ�W"#������cæ��Prl>]��1hE}.\���X�r����fB�S�Fc_	�i�#-l�0��?[3/�I$�|R�'�g!R���n���C����v�}1[d~��C	60���`�f_lU������~���G3�x�^��M֘wW{F���E60O��^��z�%����}g�v�{>=�S9�e�X�D����j�C9��_��`}>Gn�%�}����QE���? �g�y�Ǹ��st��\���e�H��>���X���Wϔ-&m��`V=����:��85� )�ԁo�┈���q���R<46ull]j������˾�#Ư�������{�dm����#�-w0T���6mcWܦͤF�[ߍx"��޳�^+��F�d�P��A�'�$����p7\�,�w�wk.������E���)[�^GL����U�^rj���Lc|_���񓊶�1|kC���b5�Ť1d��o���J��ڸ��]��CD�G��e~k_16�f��Ē�h+!�O.�>zc����>��/��T-{��s��8+��Z�ч%y  �7!��+k��^&m�C_*�	�v|�.�m�u�WۤXo�MV\�(lp/#3�;�6����G�ih����W��t�[/d�	@�GX�F�̸���~�a�[��*���y⚦@+��ͰqB�b�e>KF���ֽ�y�%�ȶ�>\��h�"��/nMzX��`�xN&��u��g�fR��9_v�6���7�G#���.4_�_u1�SB��vߏ�~����ή�-rc� ����wA V��G�H�	���H����k>�g��ǰ�X$?���o%��-kE�ʠ��cA�C$.��)#��S��n:�={Q��uG(}��L�?W/x�[(��.Xc�!J�0䠓J�lƶ�7ʢ6����&.d:�^��b�_��hZV�;'����RŠ���������D-���T�d-8{-�Nr��5��;� �x��i-"��5�=�tL�N�G^��<�(z���}�����ηz?UM�-2�v�2����`<����| ���Xe��mpW2�D|cc�3%�xFq�Ϧ�RLD��� ׸_������y��/(˜�-<?8�|!x�U>U%�ޮ��G�	N��%f�����O�@��_zI;=�E�3���t]��'
�Gx�[ă�icG�F�H���W�f�"$���S��]&p߇��
�5o�_S��9�AaB���O���nQiv�g9��n�q�LD�����P���Q[Q��Bq����W�dM?��`���c*��G44�d��^Eǰ���j7^А_��N�����b�O��ur�W+�9WP�
�i��;���-_1���
>>>�Y���G@��լ�vT�^しPn]/�A_Oc��$�$ѷV�T)O�j8{:O1�x���#"%q�oGС�1��N��ނ�����"����^��J�`$�{��u[	Fb1�5�å�*v8{��\Y"f��Ǎ� �������f����NDע�~y�qs�Ҝ��{�(^)0�n�b��g����{P/�l�F]�(����1,HE�@�A�qX���_1sߖ���Ue�����a:G�ث*��.�d�}�"�HI*�E�M�JR��؏��A�La-��������0���u>�f�2yv��J����eH�q�ld�|ϝ��:h�K����Yh�֘&�g^�f�[��	&�`���e;l�3W�C���"T������_�9�U_О��Ӱk�F���7(WW�m�ľ�J�5П�qoG|�s<eИ����M�r���C�{�B��I���N��0���76�[���cC�Pi�"���s�R���`�3�A�\�i�Ѩ�cH7o������AiN��P�Q�g��bςtG�~�.���+{'����H����҅��\c|�T�T�,�u�>Y�<��6��f���,���nBaD^O7R�o���ӷW�ˡ�q${z8����yYfw�~G#k���g?�X�h�~Ł���;a���f�,^��\(\ӳ̌]�2��A毴�=�u3���nI�2� S��*3��ݐ��1ِ'Oű�ĺMb��v�a�n���X�A}|��gf����B�����:�?�� BhΟ��~�����-�Y�W�,��U���ܼ]���<�erL}�Y�|��!u��w_2q+�;=��.-}�� r�lv}���h��^�8�@�6�= ����DY�r�~�	�(�8y���`�x0^3�h�hX�p�gg���#���'� R������&��H�F�zj�(LF���}��I��* Y�m�I	/xG�۶Wv�Qf���Z:�m�Kh|Yi�(�$
',D�6�2r����h�Dʋ��J��`�B�d�����W�Rj�<���U�sKn��6	r��2�#��A��1��%��JL�qm(D���&�y����3<=L�&�ȍI��Ni�=66x�bC�#�?Ǔ�����r�t�)x��*�p��+��P���<��]?2�A2�nr�a���XDM��C���nwE��OM�*�b�7�0q(v&j�8�],���5����[�,�W����v���/+�|(]HOQ]z+�Jjv��륛��R3�x�88�?�Lݍ�l��Tߐ9�:��P֋>^�s�����~$?B;n����}@�$ �}����$cA�|���7�m��3a�ϼ����9-}Oˊ���7��t�E׬|x н�X�'vxNo�e��)���Գ�[���6�O���$;�Yx�<���ڍ�n?r��H�+�$`��V"�m���wϭ�W���;���߳��ɫ%�vV�pY`_��?�����.��/?L�p�-��%^�"!�o�9E��s4ç��~�y"�,8A[�vDp�^�7H���Q؏����cne�,f�~�bi,J�ؤl})��	�<k�;h% Y�y�P��R�MQϠƹ�:��c�������N5��"� ,�0Xl�x��CQ�b�)Y6��qk��aZ�c��Y�H$�oȐ����$(��>:�h�p~�(v��8��ӟ��]��ػAj[pJ�yݕ�x2�)Q;K�'�|*���O��S�y �TȂ�Ioۢ��"���c��x�3�� ��`;(�Z2��t�1jLSЮp��H�$�1c	����|�,"'4�Z.=w�p��$�O��ޜ��"F!�bH�)���,��f�b�`�)q�`�����zU��g��/�%�R8��D\p78�)C�rV�!j��q���.(Ief>n�,�F
<E;N�"��ow��`��˖	Ӂ���vvA�C�v��ɮ�>oC/ًzz�lm`Lr���2��1�q@e�d��g��2���c�@�|�c���T�G��WU�(�N��#�dk0��Co�\�WT6��<*�a0����eH�LR|Y1]Ua�52��"��]����~�b��v��3t@Y�����,b���t��|q1߸�R���]�bV���S�����/e�J�Y<����G l�.�i?!�{�,�)���xs��i�F>6L�q֧�+�f.`�	�}����C/��}5�v��C�����������{�ɪ:!"v��Gi����ա ���n�AB.n^l��ǉu�-�+ �R#3��S�뱠Lv�?��ՈZ�{>Ќ��ּ�� &OX��N�Бb�U�_h
��N.P�9�l#����,��@@ ��r��DZT�`�ǡr��%�)��La�ij(��:?�����q_���]u�{��Ћҫ/A9x:�M����1�m,3k�Ri��%�3g�N�&dΕ�i�6�z��=�/�&O9�Ni���a�H'��P�$�)qХe���ܪlLZgn^��S�DS��!fk��~��vsy�`��W����7��%7�N��L�L� .�9��GT���8Bp��#UK��9�����R A���o��I���F�~S���c��Co�w�6r�u��c����m0�\�ƒqٝ�,��}��,,M���K.����U��`-���`��1��g��L�9�c�"�f<��ó¶-���m���,#��}���v�%���`e�	m�vr9T��U;���r���r��3J�z�=�HH���僓0���	>w���>'�x}_<�+*���'��n�y-����m�Q9�?B�G�������n�->U�H��-��6��Z���)�ov��m�lY퀚���r����D9f��f�ǿ=�n��Z��d˵a�����bd�}�:෧�uvl%��f��ʀ�y�m��	_gy� K��}���If�|ۈ;6�{=O���	�'E6 
�:D��l���|v�t�;��W��<M�A���A����!��:��q~��*�`�G���_qS������ߞ���KN�uq ����^�FĚZ;A��'�:\���ݾ]A�)������2�PN[��h	�PNg�F�����.���*
�%܁�(w��p]��_�}�w���?G����H�r�P��։�8�9��X���a���-7?S]�W������?L}��톞�E2�4,?�p�ܸ�X���r埻����Ga��EY$'��c��.=�x'C8	Ӓ���t��] '��I�9a���<t�4��h����Q8?��h3"`-L�2������v�A��1�1D�[�9���� c��v�&��P.H=�_��3tط�y{qnk[��ĕ�����"������w&�7o�Uډ��b˷*��BQ=q��Rr׹3s�BTc�X�w���d}e����L8�"����I���W� %�Fi����|��7�	���q충�I�G���d�d���)G���ߜ���yR{+�Z*��,�ju��KƘ�m��,���̵��V�rN���$�S+�����v��a��zq���w�t6b<s�ʪ+Yr��`*�z�-�*T{�_�*bcxiS��Ě�w]�%�o�ь%�K����7or�f��j���.G��gW���r��P.���$�k�%]AAw��9?�v�;�A��fa�*�b5�K�0��u=>�=t���!"�~�����ՀK�����#WW���լ��Dx�?�6>�tk�
��p�@C;�bN_|D��q��/<;h����I��f��}vegg7���#OQ�����:8'�0g���]]�A� �b�ymL���j��jܢ�Q�E/����dR���אt��gV;}m#�r�{ɔ?#�c��^9���FG#J)��6����1��'S�����,\h�Q��b�+�LB0.�P[cS"����^��1G��C��_���ϝ���ؐ�x2�y�AG����:`�
.~}����%�\�G��kl O��+��P��3
�V����! u�EԜg�������F��Ď'9(��!�ވ���Q�)�	�}�
��p�m��]�l�g�ի�E�O������'v���h�'�Nr�r-M�Cf͵���^��K3�|�=��_M�vQX�у��
�UA[�m���ʔ���;nW���1�T�BZ��m6[�Â���'��hܙN[��g���b��~���w�������IU	Gjo���xo��g���B��df=sɎ��{->F:�,��
��}�`�;`�^).w8˯aQ$) �R��u[2.�W[}�YY {_X�-r?����mu��G����F�E��{�J��䜷Ԋ�p�0���M3V�4D�Oطt�~����mG)��ٗc��L��	�������Z2h��$=��7���MG������wl=�#��Z���֙yU%p"L��P��L�,����_uۣa�ㅃ��I����F���!@EZiZ|N���6U!�%��7A|�8i��s��7�_�b�i�o�'�ս��s��m��ʕ/` ���^H�k۳i�;~7��5��x�L�E�j�ev鸖?���=?@sw�����ne_���[K��������	�B';��FC�\!�H��.舖�Q�v�(h�?���8�ĺ��|��ыp���9���yRҬ�� ����m4'��J�䋗#ߥd/^/L���d���EO¿���S)�u�*+E�K�[�t�l�XP#��6d�n������}ph���/B��AD �^M�Pl�#�Cw9.uQ�&0��]��!A��j���!`�QX\�9yB�	  �hrez�`T*O����Z���_��eF/�z����L�rZW�0�r,D���h s�+���)J8�2�����ʬb)d!�X<��D"�xxt�O����{�0��ߕT �*�E��xZ|�I��*y�W�`o�]O9}��$�����W�y�Bs�����i�ד\)'F�o��!��>B<@W��<255-6��{Xl���ӣ���hhh(!.~.33�9���3���B�*珊k�lI|�5;�'��O�#aE�'��z�6�:;k�?C9��,�
+-4~����Cs�L*��b��Pr���USӉK;f��w3<:���feb�Ri�j�~��,�#�[�B7�o����<ԕ0���2v���z��<hg��N�1]�%�N�Q<��dK��Co�;������D��v�[4ʕ�v!3�;�\՘���F�ꮀ�X\�:8ک��o�']V0n;��I�������o�K�>�nFZJ�էyw�-�eH�z�����T��'�����h��>��亩k������>�󊤈��e��#)7�{2<2�^��(�Q@�g``5�g�=ܪ�#��f��
rUY��H�e%�����^�~&軯����X������|E�Q=���T����~�A����˻D��)y�,�NO��pk�ތ�B޼�y����5NLJ�S�}����̣�*$���R4��p�Sr@� ��C���	������t�wvvN+��t0�� ���I�s®�:���"��BcT���1��R>��hC�U����ۛ���,�`0r��5h-����7�΋��w��;��e���?���i�x�U�q&�(+�����;�WW^�i�y,�t
�q( �-$���}z|��� w�%��PӐm��oc�u&	���A�<�# ���xۮd����x��{k�Wґ^�C�>A�}aH�o���F�_
8dh�B�W������S__��3Q�dt������pgl����k�끑0>^,���F؝߅���<���pR�I!��Ƿ|�%�s�}aL]]}�z����o�߸�o����y���<����~��wZ�߼ys�) ���ye��aww��h���A�'MMM���� ����dy��S)H`�a��R]�����6
��ӑ ��T*u뗆r��N��T�w	5��w?hx�7�������֗E��qp���,�h�9[[�R�b��<r�U����>{{{6�o�[��o��@��(5͙�h˅�(�HR�,�в��cMFFF8u{}6x�ke�B��ʋ��¢Cl���I������>�@���p�����i1*ĭ��t...�\�]{�,.j�d{k���,�ܦ'̢?qD��d�NMq�ez=�������%!��h�%�ޏ�J�0���������.�b�1�zЇ�7Iޤi�[6}Ӂ�?w������E��کr\z�40�7Po��ʵd�ɻ���]�V�x.���w�����z���rCr~������>�ɬ>/����L1C�wA����{9��4D��ub@��^:�;~�jjuԝ%�j��` ��&6�;�շ�
�u3o��<��`�;z98<�ld�e؝.+���ڛ)�0�4��6,{n�X�7,6�
�c�ư:����=����.��T�W��4���g��'���q�FY��	ZZ��!��|�Ý4���]�P�
�/[c*���~��h�8�Q�u����1������-�Ĵ���ki�3-O4�H�h���<w��^���uB��#;?u
f�7���C���%����ʿ������?l~�_6?F�����ǂI���G.zb��%�شFص�?�$H,��3M�l����e�u�%��s�5ח�|Z)�}�l�����d���矤G�F0��	�3^�k8b)����p��_�u���h
�S�\&t��;.���|,�|F_��N�P	����N���A�	S�)��GW�����tz}Sݨ�s˯a�O"'Nt�W�(�Ǘ�蹼keo	�dMP�E }�4��sSGU<�t+I�xX��Y��Uް�`�{� 3���HQȤ�j�@���ӸM9����Q�o�_A����%7�"���#��JHw7�	�9E�4�A-,W(���<t]۱�4?�l���f_4N�k��I(�c�/��U�݂��	]@�z�Io��<L9<U��!$�_����������K_U.�ć���#%��w�M�|3�t�s~���Ws�uw���z������gMحA'�l���|r�u{�9�
�����a��v����*�������X{\�p3∄2�d]�b�A��3!�FIY��C�A�@��יh-�h����U�R��,�K�:�&����������3�h�M3֗/i�j�������6s�j$Ia�7�V�6k�I�ͪ~T�?��Y���`�-�bm������-�= �0��/�Xcr�A����u�؁���y&0O�	�lǙ�����A��ac�Q���:eH����MpR&΃B����
���e�����u�/ҽ�"�}����QQ����H����D��&Z�&��E�N�i��S�w�!�y�ڪ{6ѡa���lk,���B�u7�k�� �#��e�*�F\����9o{��ߦ���MN����m��l]l��6����V�9���b�ʴ�JǶv����������cW{/ ��k,�6x��MW��D��I�@�t�8<�K_e$�ne����.�#G��C����)����gW�~�]q%�����ѱ΢�y�el�������.�Q�/������c����䌽�cL&�C�Ǟ���ԛU�,�)Y�
^~����mO�.��[��~̾��yC�m b=�_1"�B�f�%�)F��|�>���3v���%Ӭ���Z�c��2$b��1��=U�s��Z���dƜ���������]7��9��L���>�$�]�Vێ��4�@�D�]�'_���9��ŵo����옢��O'���)�����o���i����"��n��i�E���vQ(?g�!bs#VI'��{�9��&	��[wC�Yw�D������Ex.Y��,�]v}͂��3�F���|HJ�,���zĳ��F�3M$\���Ȣ��h����O%陫�*�.˹P�n��s���B�%�M���5�t���|�^�s�t	{sY�/S'��2� iI�a�/������=#�#<!���%=?u"�n[�b��E^�y��c�5W�<BX���QL\��IMW$��4�5�陀��)�.H��|����0�@�ɐd.~\\���/,\�t���P��|�6��Ѧ��Wd����a-_�冺:އ�(�QH�n%<Z�r
�9b��㏞�!��0�Qz6�C������>no�nI����+@#����5چ(@j*�~qk8���?�{�o^6�ȓ$��\?��3�4U����P��o�"�8�����������m�$��J#@ޢWK$��r�	AFʝ�:C2R���E��}~и�%a�}Ğt�]�$
b��Si��Տ5��N�q�qf>
����lW�
e���*�>12Ȋ����c�& &B�^hз�M�RI=	5�������[L�Q�m�K���j��Y�� �a�u!&ц^Ae(5O��v�d��5��!��c��e��ӽ�gg�N�>�Y�:j����g�>�>�&Jtѱ(�C^8�55�'���l�m�.چC�,9���N�:�'�=h���D��`}�,�wSh}ᇢ����~�܈�}�_y�N���[����kN}Ṽ�\�B۴��OM��g��k�d�-9z��_8=��^�G��M��-O��m{Z���Z! ���,E^�/j��`���c���϶ěH5\U�LN��h�40�`A1��nI������4ې��-m���x�:jD���3�[���
)8���3K�cl_��L�L���`-��^D�ho�Kq�HM֏�F/���tO��=k����N#K�`I��=�p�8gV�Z�/ɘ�#��PB2�G�e��HۄW��v�a*y�!3�V+�Z��p�6	�b����\�}djaƷ�d��Z�CͶ��̤��W�h`�C���W�PZ�T5S9�\ �o���J���t�Jz��H��������Mw*�}�)�$Ⴕ���Ԑ�������yO���S��� �7knA���6h*�p�!,��4�[�K�c�B�w�<�\�$���V�Ee%�,��&t��t����_�=z�&��i�R	�έz�����������ݴ}���]<Ezw:^Q����	�N���m�y�
� ��� }�N+
3�@(��4���C?q�rb�/W��b��q��ՊA�9"'"m�h������t�	#�s.ͥ)}��6��ٽ���. ���5t�5a]��oNE>�pY�d��	O\�r���\�<��ݴ4�0Lc:���Thv��u�����wdٷ��sz//!�~�Oo;P���.�i�B�)����@���������N��������n:xL�!�F���ӭ�(�O6b3G��Q��O6������k${vꁽ��I��y?C^�l��w�����%(�t��{��F�Z��d̪s����jD� ����yw+��Ƀ�_�Q�i��X�@�M�t;���~��(������/�9�z$�¬A��ө�s:�K������k7����m��H��?rĨ��R����9fk�L��\C_�m�E�gDn@z��`Q}qdo������� �|�! F>�*|�L��a 5gk��N��ī�!K�������:��+@�O��?��H���!xvzmj�'��#�w��v5!v���dgSW���}�L}Jؒ����kT��v��w����(�}��D�oT�g�oHS�.���h6���hc�v�t�#�V`?4�g�@l�z�k�
�Z���H���_C��)�LGn�f�� C���p~ͨ��׋��\G��!�.��HI�6�,��d+��W�`
�:���E�x�}F]��6Y�dE����"���R�P��4Z���)~�,�3���u���Y��s��
JLԏ_D�.���i�~�`1U���k�Ƣ��px_��{���a���-�u��\�f����*�O07���*}�s�l�Ow���60�)~�Kx��^����j��1�K�1�o��񷁀>$>�}iz�M��Җ&�ٸ�I�z��]p��c�p�o䯔d���e�}�Fx�Τ|73��=��!C�Z��$|�|�zތ5:k����ֲA�8�Gd�k�����^&)�X�&���dy����R�����_��$�ۜ���iMQ����l�ح���N�����������S��7�Ɓ��uP���9'7d����;{��8L<B]'ĵ{��}����zbr�"y��56��a�!lY����O��9�g�������y��!��n�o�)��?P���*py��H�^����D��D_=;���YR����f@��M�&���wVcKi�H��6e�V�/�΀�����n:��8��F-�o$��)����{ٱ��\���ۋZ�TQ$�0��t&�8ٴ=�G����zDӖ��R3���,UJ)x?��oB\����ڽ���v͛����v&# �8��o
�,�o�N�	$��+[p��&#ϭ�>�m��E����E��Jk�p)�lK%�^U����Hb<~=o���p�� z�h�<8�GR#��w��ހL�u��1����~��W.��W���h����kz]p����`O�eM㏱Z+�꟤���;�4�%\Y�m@�ϝ��j߹�������[�P���9ٽ"b���a�'Ϋ�����g��QJ�>Ә��҄��Ls�������g�j��Sb�)���� &�,/!�6M&-�D��b����%My�v�7�y�f!W�&�A/�<�5q�]k���dq+������U�k�ݣh�"�V�V�'���_����q,�y˼C��V<���\}�g��#b���\�ܠ��÷ѕ��tQ�n���W���V�������z.A�ٝ!C�e�J0��	��[MH+ہ��q.�>}�\�^dY'���g�,��6L��T�a7��S�z�nO���XǛ��f�G�9t+�F�z�F�4�~���=49�Y~R̴�`��e�<��I �zo�i9BQ���:ٟ�'����vp<��;�?*��kkVd���x�`W��/"B�*u���f����ޮ��@���<A{w��4"_N�ծf�>h�˾i���<�ؤCf!�<����:w,j"}'����������$���*�M���#��_�4��ejNq�p�>��.&`x����|^:Yʗ��*A!j��ޝef����ݦ��!��Ds��9J6��[k��&d3��F�J5G.XMV���M�G�24�X�"	��!��q���3A�ʣ�q��e��Gق�c4���H�R��l���Nv��n�e�S�l~��3^Bm�{��i��n5
���x5���w(.��K��bsǒY��=[�:���y}b��7�0�܃�p�	�����Di��ׯ�nyC�XP������0CJ�])�C�9T���cS�q�hЍ3]�)%�P�QcF MV�'�Y "�A.�G���~��r"��Bd��"���oׯ@��D�����-v8=�qqQD���حH�d��B5pT�}��[�L���Zz�Tүy��foh0<tU��5#������XzX�.�ǤN��R�)����s�>�Ŀm��8���ܭx�r@���N���?mȿc�Y�J�����iI�`�����e�Yˮ�uS�(�/��#�ua�=���{��H�H�H�a;ߡ�kv��NV��Vhj��>�������۪7q��}L�_��)=_Yj[�F�ҡ�}�B}�K�(L��o�T�t�=1�y�0����Wg�|v���+��<yV˙�F_��h��U�n~��5#�eu�b~=�V�vYW�I/ȅ��!|;:��{�xW�t��nɱp����w�j=���>yk�[�EY>�ڿn[0���<�����B��k�0_�P�����E��Gl�Ql��خ4���B;~��WU`�����CA��zB1�Lo��H	@���-��s\6uFZ����
��Eܟ�C�������*[�uPI�l1(�B�lY�H�N3�d�H��![��(��dc7�c�����~>���q�����9��/��q�%	���]�	Lف���F�<�ן�Ƚ�+���4e�6I����'e�eܹ��h��Kd��?��ț�Z���D�Y?j�^�(S��q�:�?�i�q�	��]����J��/�Z2��	�
�@�(2g��h�Ԇ��U;�~e�-Z�{N֏���?�������7i�5MC�>��.J1�i,0�Tew�=`[�m���tt�w��I�E�H��~B��>��x�e�qAC�����i>:æ��8��nK3AC���Yal�G����̓]udn;�.��^J���;`�����D�bZ�?� 2�9=,/4���(�g������	<���]6�U,�L�@᲋��I�)�#{Y$��Z��ˇ`zq�(��t^��+t����p�	����gϵ�}�,����L����Rڰ{[�m�}�Mū�����gg8h�Ae�3�[w������\���� `
.\RTd�R��e-S�^���/$�u��P�s*{/_��[]�[HS��XnR ��V�"�d^,����hs؆R6@+���)�W4�����cI�{���IF[Y��+ʶf+�A㹐W�uϗ}oF���cYt�hͅ:�uKB̴��9[��d>�4>�4����P8�Se���S�6���IA���Qh��ۻn�`��&ԥW�9k�a�'v/�{��������;���u�X<@�=c5N��Z�g�&�*#?@y� T������Mc���I�$s�x�Jf���	���$�}���2�׈{vΒ%%O*|\.�L�T�%�iG/��z?�`&���GE�DU��O�[���$�k�f��;Y�w���:t���6�e]�bEj6�����5�{���+����P��RB^^�����'��̊�&�6xf��������W�8�{j�	��2^�A%�y�����H�;���v�����m�`E]"��uc9֊��?�8�?��5��i���|U`�hh�=��,wﲋ
�v�^�5�;K�-,�PB�>�TXo����u+��S�zUZ�����t�L!�v�y���L
P��*r�&˯z��JE�@_�ox����p�ٿ��o߬ %<��x��h��_Q����Um�����md9��B�_0�/QqéC���LS��ż��c���Я���C����i�����B.�K-VAۯ��v�
�w(n�����F=ǰ�2���@Gr����Q08eA������w������mыs�	߃zZk0�N����"��+�-84rFİQ-Nd���� }H%"�5[�\�}a��x����0&!V���q.,��&q�]�S�<�H01H9�ճ�g��zfh���k2�WOM��ۼt%�tBk6��2��%���x��C0Λ��`u��t8*Jenۉ+*����rgi>�'�kT����z��;���w,d�H�pxAr��@6u~	`¾���Us�S � .�k[�=ϴ�a�c�O�/��e�5Y�G�;�D�[���z�� ��Q�/�2�R��Z�^�r�U�9��������G�~淲&�{#�������Ke�^��g�#� �ܐ�9���t��?��N�J���.˶�ZI첻�)��!��`RYU��<�8EW[
0��/j���H�&��4_��������Z��	� �P��-D�Wٽ�'M�ћ&��Tg�\����x�Nż@��i��mD,��N�)����%%��۩VD�&D�YYuT~��^˕�3\���M��������C����cZ�W�¬����!��T�9h1�U뜒�g�C�{nz���~�Pm%�Ⱥ�z���������|_���M-\����������`�{���XK��R�?"�pƲr%,�Ŕoy��ﱚ����10��nն�v0�E��#^ �-
�=�b�2O/LZ�Q�߸t��Y��\/��� �|�L�D ����{g����;�}�-Q~�f�`�n��Q��Er���cuj���-d�g��g���!kRq!2{��R��ɛ��S5�s{����'.�W�6�|��(�����λ�w(_��BPU�}�?Gw�{Y�����~gH3�
e���}��O�j�Ʊ���t�q}*�R�|�N�OU�&�Z���E֋y�o@��|�h*����)�֥pB�wF�y�\l��bL}�rM=�e��$~��q�ao*e#�4)f��o�A�&�5�)C�a��iWwש \�Fa!##C�%7/����D�L@�F;��h�5��������~fNfH^�nt8G�C��-D�>^3�&�,������$���8
����U�S�Z߾�~�df��B�x7�e"���fgǆ���]E����������m�K��ɔ�\�C�5����tr���n�N��o��B�����ĸ"AP9�B�S j�N7��c���J\~;�ZS"��9��^I�O��v�n7���,���52����ʰ�i5e3Kɺ�z�*{�v��sB<�b��yƩ錙�����B�V"���4�3��܊J8H���t�7����s���	�1�����~�N�^�F;��/F�9鼵27w�2�S��}���ȧR�ഷ����l�+���سZ7o�
h,�O�l�qq�Zl���&�
;'Nnc�z�BPvi��;�.񪂡�D��(�����=4���k2"�>��o`WC0�]��(� l����J:?��o��3�����C�~;&U�S^M�J�T�NB}"�ǃ�4AA�w���w{�3zظ4uF��`�����?��5��o,$ay�w�nc&f�(�)9;}�����El���9�"�/���>߲*Qug]eW�	�f-�pReo',VRrD����Ũ�&�kr�x�)���mMJ*�G���h�ݯD�`o����t��]����w���ďE�+L��r��u�b���{Sđɼ�Y��y���77A�p���}0����G��!s�d��p���V�5NOu�V�?_t��M�����,��/��V�S�O�)�,��yXE��:5��~!��v1��+[�L����=m�$o�!F?�	�����}U`�2z�--O�C������t��L7�3��������b[��Ʂ��~k�O�Y�JW��9i�5�$��>��xVA_x�q8(o���nQr(+���T��PE+GN~�ay��B�)�*C���r�A?�P��7̫R(�Z�1>1��g([8��u����Iy�C�����b?�f���ҲD��}���/:2i'2��
�I�n"W���!J�]gpc�;�<Xe�}�l[f�-5�y)̾Y�ߴ|VI�����Y�"~.g��\����U��M/�:\SN��8�n���lr�:��;��5L�?�DY<؃��S2ӌ��Z�	l�޿��e�عMT�T\�[�M,��sAٷ��	#��W��l�� %Bc@g@��ZM�j�.T��[����/�3Y���f��B2��B��M����E��W�4��d��x=�����j�)��Y{�ޜ��1��J-.���Ji�o�z�K���fX�Q�?�3�;+N�`�E��<}�0h��Ҍ�g����E�Isa94�V�C]�ep��q�a<�	F;��c�����D]g_࿺3�hʨ�=�,�Ҧ�,�(��?x�[\���iۅR3�祏���B`�.����xڄZ�+,i�jV0���O����D]�V�ˣT���:�ۭ��Fb�A$��D~^����Q~�u+b|%���t�Z5"����c��*�����.�RH��G"cHokw���3h�S�Tb8���#���+`�@�
��&F��,^��w���dI���}���W9;Q5�q���5��u�6)EK�/�5�ҿܢ�M<��`��[��.JiQ�0����ɝ>��ߊ���ސ"7�Y���#u*+���U)^����ຐ��7�8��q�z3�u�QzB6Y�fBb������ �?;ښO�m{[�
���9��Lu�����~΄��Q�<�r]�+gA%�KBG�@��.��]W������ʉ���P����T~� K^�`����ݧ���c]]%bV���i�c$��	W.$�zfStU���U�9�^�f��᫕#xl�RZ��SY���A�����M�F�� �1��oO�{�����VQ�S�_�9�ҏ�eC7��;�FFM:|q��U#�*`����5g��l�5k��re��=�ma=�8���2���{�	���2�Fc�e鳚����r�gp�o�Q�~c�UI���kWe5ް��Y�j�᦮vZ��b��>//����+!G���|
8A���/_x��?�Q�`E�������ߥ�#X`�
������ou�*}��"�<5��6�#��W�qf��*ߐjg�j�j��s�F<3d��9��O�9��3��lz�ҚD���T�"�#��R�g�W�69�v���������<�t���1n��լ{����}I�T�P(B���dz�0LU:%�]9gԬ͖-88��Ƣ���a���-㕘�IK�����4�>9�3F��j��I�l��K͕�|���&�����ᆮ ��1�cNßQ"��`��{�$xoR��(�F���oLi���� � ��Bp浒lU�
���K����I���C�vv��X�^Ո�eE��oe˪�W��������%�_�*H?���~{A�<��r-���`u��/�y�rॏ��6�K��L�U��掮Zܶ*<�(nM�9�-��gA�/{���.C���-�����m��C"-W��S�(	P������[&�-����'�V^�nd&�.F����P�Sm�-Ql0�	5�A��a���[!cصT�{�e9���oё��N�W��B�j��K�F )]��z�3�OI8��j���OF���}�S�(��π�K�iX����1+����ȱ��k0t���]���@�i��&�Q�C)규��X�������(ų9Y'p�>�Z�Eb{X`�w��4E ���)��硹��izG���Yz��$I$%��q�ú́hA���{�ŷ����~���/���W���P��~B��u��@Lu@�e> -��+����A��
%�,�K|iB�����!�+��w_�z3=���kN!��4g)�q78�i�ŅS�y�������P�=n�������@4�)VZ�v��VK>_
��g�]AJ�����Mܐh�J��)�h�����lQ�ko�����ύ�����>���BEd��]�H�
g��rz`��7B:Ac�=sw�����VW�<%br�#+y�|*��l�k[��;\��pvX�"��1�u[���� قCvj��=}Pjv)�#�nAF�
��WI	v��V��^�atc��`�����_��|�v��:W���?��	���t?��Q�z�
�\ݸ��o�bG	� �m�k���"`~�������E:ަ{i6V%M�鳴�k��'�w0��g|����/�"D���U<x�BAc�ٍ����F�s��7tV&���������Q��2�F�����R�ڞ��mc6�zu�Ei�W�-��D��3��,�3k2��{Rd����������TW�rgbAl������3>��5k�-<7�<���U�q}�oKy�֎�Hr��J�?0�	3ܡ�r,]��8�BVoXf��dy�\�UZ��o��~u���U��Qr�!E�}=}8 -�[Z��6�;-�T��v�����ul�vUH���P��2,���p_��Xen4�[Q��/<%�ڰ-%v���<�3zπ�wTqka��i릔���>x$ήX�К��r�c�B��*S������a��?"V�l��4�ӗfc�?_~�V�%"R�'�����Ң}{�(��a.q�m�g�Wk�KQ:B��6xs���B���#S���~�Ns�9'I��rE��kmV�݃�J�6]*n�DX��\�f���tY�=��Y!�Я��_���MK�S�Tfæ��~�^Y�b����^�G�8��ؘE��BH�;������p&�/��� �1{�f��5}ލ��!��O�q��H��h��q�ZU�n��~B2%g�zc��z�˷��gx��o�|��]EB�p)�T�.8�����p��2l$ ����o�L��g-����~�k�/����0%��I�finn�|4��xh���'Sa9�u�m�r�3��f��g�\B��TT��&�p*��-��\�ԓ��w�a�\���m����66Q�r) K7?Q�����ۀ{kf����cF6Y�L��|9����m�C#��D��v���y�)@Q)��܅��k�e����_����?u#�R�0���r�n�9^��j�9�VYR��5��:�q����w��}+��&�s'{��G`�th��z��dD0Ȼ5=8�b���1�?��멎aqKF]�$NJݯ�3���j	�)��F#�t�����4���,�	�rC��3��+����@ٓ@!r�{�bٶ��c���<��0,�4��J!�q2��{�	�.��ך>{�6�L���]o���d�S��^�����a���@ЄP��	4��xO���U1����J�;���u7o6�z��G����������)|H!���TxK�����^>C�R�����0���\��d��\��륥l�Y�k��9`�z�tjP�;�3��bY��3߃=̀ή4��蕬>�=�M#�΢��$O��`�bs������l qT쯇Q�R�����%�;]*��,���~8���\��4_��S�W����Q}��c
whLea��f`�;>*���0��l4K늆�t4�F^JG�����P�x4��W�:�9��7��ӌ��Ӯ�,#"���0��ɧ��k���(�4��=���ð��Al@��b�����dGY__e#>(���y����	=U���G���4�!f���^f��g�1L�<F#��xMl?���"�*��G:�^p�����db� ��r�T���)��|qKL�6n9�q��BG�5�µ��|��]H�C�?s
	�؆���O��̎��	�c.<������(��d㺑A�8p�]5�!��h������t� ϛ�Q��g�|Q��͙z��*����i�&ǧa�1��չ�W��|q�FL$�:����~�?�U!������)�����,�@#:�c�����ү�O`�[����z�溂6}�43�Y�+���s
W]�#�.����F��*�����6��zѦ��#�t:!��D>��6��&zCBF	e��ne�\�~>S�^AM�\����l��p:�tNbTq�J ��Р�}r3	���3�|����C�܈ �n$�	x݀
�a�J@��$��oYF��ɶF~_w����Q6KE����;�f�ۜ��=�L�NY"�@L�#��fð>�=�Q�z�`��x='@��B�t� �(^1gm���b��C�OT)�my�Q���Z�Uݨp�.�9��t�d	s}O���}i {x��V���ңp�;�q*�XG�S�U�<��PƳ���=���-�s�ꔷ�7�GM���a'�@MN#B����䷤E�Ɵ>j��)�S��9F_�q�O�3�G��!�~�!c�UܡAf��&�^RຟqM�g��c��$Iƿ��&���5h:��ڱx394�cP>��w��ӛd_��K�a1����J�1Ǵ�$�#�4��<��A?M!���)؆�	��̼��6���
�He74&��M+��%|�kfE��b麀|���3��A���ۚ�����<��q�n�Kt?��͆���:.
h�izT����q��r*T���t܎�"q��_g�j�(%oq�r[�$6��M�`�(:�9�"�@a��a��k<�ճ�2�ԦANP�����E��{�>+���g�vV����KS�w�p���fh9�8�u{����-�%=e揥�\+ҍTe@h
ʻh�MG<�oz®�v�.jֈ��{ϣ���s�-���f����SH��9�L�G�c	E�:�>���|�?�ܞ��n�g픤Hgy`j�MC�|��y���f/�۱mb6��8��~�3�������c��a��D��.$l(��D�Ҿ7��6�����g�@��/���֚I�Μ_��O#�#@��%<��P�<Bw��i~R�c�"[%e?hVi�=yTOQ�� ��9xF<�xV�9�}rs�Ú��'I`��oKQٺ�"{��UVw�T�� h��� �h����<�d��š�[��Z�����k��9��+T�*?��h ��n��#���������۞">��Ђ�� P ��2xD��"w�jw�!�c��v�H��{�)=H �i��*<�e���ؓ&ǘ����c�����;�����,{yC0��37q�P��u���W���k51�0�v�j�C=�i����nd�w��;A���{��}�.�v��e���u{�&Xf�d䃰n2����i��v�� �ȡ+M/��`�8X� ��b1�`�t���=7ɟ�ʢ��Z��.u<�y:}�
�ˠ҈�_�A�2�ȍ�|��L����,�-wm�q8�\�n��L��˻�'�\�C�^�<��;���⋋_�����nP�Aw. ���
ı�H��|�{����P�c�Z3��x�lu ��u��x�F�����	-�<�I�$w	�%՚B�BT�ռ����/���4Vhe���BJ�b�]�
��|����<�)�`&{�x&��7��[��n>�`8:DƁ�ˍ�����N�� ����㍕�Qr��A;Q��S  Va\�
�{L��z�������ȶ��1�?���Td!By4�<�����?ǩS�ǋ>�]��#}*��9�T�aA�Rp�ךj���u�ƍrW�OI^<�1EH;��M�O�u����RU��s�s6�^pG�p�y9�G��E_k(����!	f4Y�
��مtN!6A���~��x�g@���h���M��������Hޗ�*a�GV��)�vi��������h�㨡7�l)�!73v���]�7��hAll�?_fl��;Ͷ�`��5X��1-Y3���R �@�u c�@���V�"�����NɆ=�d��IckO �ȜQͯ�b(���|�}W�k""���A�p�6vT��~8�����/Q�7�~D��n�gK�0��a�?d�(qB�*�<Fq��L������7��]Hb��� ;����N!�J?�h�]>��8�bl9#�c2������	[��>8�xH��+߹R/�u�?f�|��G|��E����LM�F�F�]�(_���|gx,�t&�t��!��(^4��|!4Y�
�<W��cq<��2I46N� �k���΅�L146����-62�x��V��>I���|�\E��71��;>.���3�2�|���!͈�DASL(О@%z AA���B���M�Y��
�J_�Yq�9 ��ۅ����hg.X�4�������/p]٬��w�$�l�m�&���k

�Ͻٲ�|��,�2��Z*i
�}dHǎp#2� ����������n��S9�F��o�.6>
9~��b}��{Dc�a&���*0�6-�zJ��V�NoM6��Q�3���1���/�Jvv�O�a5q��ئ.$�2��J���	 T8��$b���Ȣ�s�B}��1Q��2�v
�%�ۦ5d!�U7E(/��0k��ɧW,�8�`ͮb������.�!O6D);Z�vh�KGz�ՍĎ�F��|�(��R��cRFf'>ĬW_2Ш2�1ݾ�2XB�
���&kV����<����Y+aX~��w{>pr����@�E�y��Jq�@�)aG88đe.�H���ք8*&��Htb�38�^��<&��"���V�b3H$��1���X�״�ү_/�V7�iO�tX�����&���C�,&�������wSr�\�t��T��[�F�t!+��,��ƴE��0�RHТ����n���2���4�gZ5���I'��b������QF�1�^��@�]3�p�$�oׅDP�Ps�b ��!�p� �b*1��8g�$�o��WG@g�7oY�9O�f�:`��Z-ǐS�E�eCG��C?�����_������Ǽ�č�8�vvCT��y���
��Bdy�j
�f@c�I����В�rM��0�����c��w�Tf�	�d�nH��h?YO�y�dشj�df�Af�j�V#���D ��<��Oc�f~>�YI����3���<T�۰b哜�� j�0O�n��WD�4�)��~e�fӞ^~_��� jt����&T�E��)!��px��fa4֒jƎ����7eʉ�"����
߾��r:��|�쟁��a1g��IJ�o���n�n�A�H�&g'֛'+"X�n����:.|��˝��U��Z�i��r�d�VNM�:�/�DW鼵� ��h�rt�8ȗ�5S���|�>�3�h/�Ʀ�>��ǧ�[��~�̰)�̰x��ܵEЪr�r�w��q�h'g���\yTl�&S��)���s�D�������D�/N�r�ͼ8K[���'�t��������%�
�ؘ˙\�h2��y�څUu����֫�W�J�c9�׍�N%n��$�O6�6*r�Sn$�[$q�rLh!�P\�nX�L�����R�����eY_�(	L|�! r׀.�:��fX+�8��+,��Dc1��C��H2��BT-��0�h␑X�W�W�)�U?Gg[��ɳȮ�G}PH��w����Vb�j<&��~�jMY��XS�/I!�4����:��h�"?4�E������b
�\�c3�W�oǩ7z��ӹr�z��7�$Ӏ=�0�K>�P��6�@�[b���d_�ř_3�^��q����l�`X֔F,��}�%���:�
:
�����%���&�\�T��ć������t07���˳�EKr�ή��QC_� Y�������(�ui��q�u�fRSΪ>���?"��|!�5��EuJ��mQeg����K�s o�l��&kʄ�Ǚ��qvQ;)�x�d�uAVs|ܘ�Hŏ�y9u!�f�ʋ��+�W� ��B(a���A�
�W�+<1�Z���/(�a o�Z:8_wB�E-7�jf��7Co �[۫�4���Ś�ˀ(��&.GW�
k
j=A��,�Q����;qj����Bٳ�mm�vz �T�����Y"�΢�f2�MN�I?F|zVOUv��}�|�	F�s*��9��c�_@�rL��`�N���� �gKh�Ǯ�N;Z�*nP������Q�l�w��`@9��V��K���b�1�w
h��D�����X2���Nj �ł��Z�~-�����n�@��~�HM�X��B����飍�H`��#�B��������v ;|a3*����s �I�dt3�|�;��{���s��"�.[������^�>�i*�k��`����**I>�2��CIU�V�4�A�A^D�:�e >/Z�n�,���T��E8 C?����Bo����Mj\2hG4�5�g^�����8���Mq��]�io�2C8DH��ԡyA���>��h)H�y�Ī�G�}JJ�����̮�s��N�ƫӛ�C*�#�kGI��~ջ�I�=�^V�R��~J��T�b*�p�j\
1��E;�kO����Ӫ���qv���ԭ/���keY�Rڑ���@��Z�5q��짢�:��붨Ѯ�_/B��K��8�?���)�h@$�2�W�����`@\�U�.�L�
�Ͱ��<�^�b{�˅ޫ�}��Uvg�rz��6��k�~�"��J��&_�39z+-��`q�Di5\��#)�(;Қ��$�.����e�v{U�Z��������V8�5���4ݣ���P��D��&	�aK����H���Ҡ�+%Eh߶��-�{�� Z�I��
Pp5b��+� �}4�Ƚ�g_CC�|��S�d_�����K*�)*Y�;�.�,D !�v��@^��2mU��5��"��E��ޫK4*���U>Fж��lh�7��w�%΢c]��+h,�b��0l\?��+T�=��xPWX�[��1i��qvXq�9�^����Y0�e`ZZ{�ٛ��>J.�qu��j:�_�:��D���b¬�,�dR��㡓h�(�E8�^ ��NK�`q��� �r@�%��=����@�|7wy|��sX�X��I�J4��CϡCW(fZZOm��nC5��T��#%8�����@fu��C�i�j��? �"n�BJ!n��,�����4��O�ڭ�D�Q����+��b�ֲ�D]>�-�Ug�Pv�mޘm\��{N�@��s�#�訞A��� - N�Q��=�e��Y�l�n�┿:�/Es�mt,d�f��@��8W�Yш��5�~���Ӎ�w-���A�4�H޵�ݍ�����Y�nЇ��~�{���8ٰԕ8eFک�;��_;q�-ִH<.��La����H<w'���,{�8�/H�q�!pD�ñs^�s�R�O���Q[���j��x�/�����C���X<���m�=��	g�ƃN{r��ܽ
��''מ޹%�W6#BJ��X#]��������'O�8#\��=�N��"{FT#����S�B?~�7j ���P�|�p�9��9��0l�r��|s	aa�aٿ�k�ڍ�P�B�~+􆪴���&� �+����Ys����^K������eы����:;��./@jOP��؁^�4���)l�q�K�2���Dٕܩ��y���.�l�]�|U��f��v��O��x�?�HA�5�����0
Il���]��ʛW(:��Tʠ��L��Q��ŧ�3�If��̊ۗg�F�Ad})��F��^�n\�Zd\��t�94��@]H=4d4$�"��ٓ�ˊ0��++���v(�N���[�U���:�X���Xg�aRoOϩn`{���E�o]���QP���e���&��6&#������oQ�FZؕ'�#�2/qE�ea��	�<K5�(?�no��@��ҷ�rD9f�+�S��܅<	�	�T�Uq�����Jca��B<e���-�	��9�ݳ՚GԌ�.�S=wV+�.��P�q8�����dbotfI�֢7�杀m0��������a|?@i��,SG��Gy�
?!���Ry>{�]=�25���e���b6#�I���bf7r�,3�u��֒)��ry�.���6~BnLO`D��tM����]��a���n7�58�-��op5x^�@0�4Hʿ����k�5��$�����c�.��a>�L�����,�4^6�繬��밢��
���K�M����ʔ��9�gT�]U��E�Ch����Eh5�;%?���.��꟣B��{ό��F8_��D_���X}������+�RVa��٠	<��	�p�*ɠY�,ꢈ����,#�{Mj���{|.��� �#�r����/v�xT��EG�:�T��X*�UTh��T5��ꐘ.��X.DP|��s�+�_�.G��pQ�.�`��ϒ<�t>���]�5��s`�����z��V\�<�,�7:,ퟐL���m� �W:8!�? x�0��/��,����!�"�,p�������v�5_3(0)�_���S;�'� qk"T��N#t#�o�뤁�!�Q�.���k>q#�cw��L9��11��n�O>h&��nYZ����{���l�Y������Zݫ�s
	!X!M܄!U��|�#���J#*\��ګg_��vJ�,R����S(긘s��b��V9��w$�}J�d���m��B�旔�� ( 4 GE��c��I���C��΋w⠗�������p&O�G�b9�tAa��G}���9�O��@ iB{\��X<���}Rn�}m3���ڨ��|��⽹���H<�A�Z�q�V�%y!{���HS�V���n������s#�'��5��W��dbe�>Fp_p@���]��,egIQa�$/����� �Q]�f�,��)]�} ��u�i �i eDM+Hi�L|����b��\4V���:twĥeP�@��2컋��JIdt��r~|���'����յ��+t7!HU*(��P�7.�Yv��%�5�)�,}�z$&E�x�KH�����P��C��+#{k D��{g#\�X�]y�*��XH���}"��&�q�&�F�Yj^�46�KC�{�T;T(b�~e�r���\�c�^~���N�(;�H
�.x���πNcK���.B�S!�ᔠ��?S��$3�p���t�������ie6��m�2�f�E����믖�(W�����3�� PT?0'#Z��� ��Y��3�@�q�����=+}߷�U��7�	�j�}�aM-�>l�'!�g��s~|V��	�,��D��gA���Úw���bu5p��A�?�:�ǭ�7he�= ��93�%L6������Nl+W��#�m�T%I4KFQ_Sl���a��]�q��Qd�D���.dY��3����r����͎]�؍,�9��<��-2�`�α�.�M�kv���նre<��ܽ��ϖan�6����j�����H��n�����
����r�ST @��`X�W�[�\��-�n���T|w(��d:�kٽ��<�T���.���W3U޶�4-��t��.��?�[����m�V���ru\F*��Qׇ���n=?�����{����fTj��+�����9U�X�[\����D$=�?�@˓��V�������4M~k��R�VS{��U�䗥�*GQ�?��9��A��<�aM���/X�{���!iMmձK���-l����C�/��V� ��jfW�{�moϭ J�؂��1��S����4���_��+{V�$9�?}�L���@�gf��p��x����J��\�p��^�����������>8�v�@K���7��֍J���4f?{�\��~��n���{�WtEb��y�;;d\�w�!r���~)��Bh�H�i�D;�/�^ S���5��lM>�JR����
����78��i�Dju���G&�CrY/�Yh*)m�ݟ�i�-�)����������6�3/����2���=(�t\tظ��4�sjXѸDd�����J 4����t)*�9���H�HݿF	��P�iF�;���h�{��((�����m��K_J?�~wҰ!{�K���-t�KH������d�Rv��3������N֕�ʶN�WU���w�b�����F^*��$�ĝpiZ���ʹ����t�*~��L�ry��W/֊[�Qm��7�0�ǟ>�m�4-�?�Y�=O����vr�B�J���+2�&�!z��l2q�����HVpI:��� a�_N���k�{{�|��}1v��a!�#��W�@_�9������Ȼ���q�����8��k�N�s[�<'��4�R�(v9 u��\C��*U)U�$��}*}Z���5���|�Źe�ϗ<50t��O��1�����8S���i��^���S�؛�u�i�C�1b3�R�= s���}�=�G�i{ �a����ؕ���@��@w�*6i��̣��K��;!�[���G��L3֑#G�����<Jz�ǂȨ������U�ЇȪ�Z��<� ���~�jlA�.M�����}_k�f/���R���C~��A~�ߎ��(ܿ�a�Ũ������(�ľj���ȶ�q�.�5��/@d�������!�ލ)0i����֝���ˈ<9:5|�y�sU�9�Ίa����Ԅ��s^L�T��t{�TY�<]�h,��/f}�t���-�
=�[]����z	��z�wԜ��\��\�!�\:p�`8,�=觝�u����k�Lch�OuN9�'θ��@��7�Er�GU�u���.����7q�3#�V��w���_�*�T?�c���z�o ����6����k�]������O}�Ɂ-�8�e*H� ����z��"	Ҽ��>H�o@����?do "��7���@r�Z��ܼ�,�mՙ�7��:��zJ�
�v�$'����';�:$>�E���q�`�nO��w���8Z��	����B5~~)^Z[�z�R?��`�44(�K�",��ƃx��I%�2A��X�i'm�1[d7���Ѩ�åm0�T7�̈́�e/,*������u��ta=7pis
'"����=��Q�f?i3\�2��	��#�|_����'T2h�J��7�����7t���i��2�u��qIiը�-s�p��y������ɓ���� �<�~��>�W��b|�"�<!2v�U;���
˫�--�F�Ӗ����u���|/^������J7*l<�W�_6^��]B�4��)ݴ}�F��T\D>a�af(x�߀ʩ��������BRa��`�_�!��g?UI:��C�i{�2�ԟ��1�߂�<��]��ǯ���y����o-�)�С�q;���9�[c��Ο~�+�6?���?׃���~�:.�g�g�`5������;?�,�����-QN�87�8yR��+v	�F�+���s.,�k.(�[D���{�><<�MdOG���DN��|���1<ǹI�Qta?�f�clJ�Qo֊1P�xpͤ4����VD�_��8<R�S�8�</��0jOKz�j����v���`�ıko�ƻ�NnP�L�0��	������an�b
dY��Laؽ��z|�Y�M�')܂�)�y�b�'G��e���)�5��t�i�AA��or����7�Ɔ���su��π6$=�����NG��`����$��f}uϏ������A�=\�����a��y������r�h�4%l���'�Ã�s�WʏJVi_�9�V�({�#��O�w�76����W�ڷ�3�9y�B]���x����\#OR��;���?�8���l]H+�������n��F������ږ�Qz� �0%h2��,憺��O3�ӝ�����k}gp��`���%��O�K�s�]'t?����r%��������T�a?h�eMr���=%�u���G�s~���t�tP��]�P��.5���_x^���*P�?�T�q*�����7(f��N�P��<�p��{�v¿:�WX�n�P��|L�F��z�a)��;½cS2J�x��N(@���6�ApZ�;hKa8>�,����)�����*7~������
#n���<>C�j'����6K�P�:��������; �I�Jc�?����F%�`��ئ#�S�!��j��!`�WD6��w-N���R� ����7������G�wmH�"I�T������kY���&{v�0����;!�ƾ���}���������c��s�Y�����7���"��Ү�'C<S���qw]y�~��_t?���%��Y�9��5��M`�bX�S��K�U�Q�6Y:N���@� �R�	���bm<qO!�/� u�#��*I��@��444�;�6���;*d��ט VU[DR�L(Nff�Lȼ�D�i�����*ڏ^�'�����������n�ь�M5A��L���v��-����s|�5S�Šh���@V����^�F�6����8.w?d��Ɓ��u��;�ie�ٗ'N~����+v���Ҷ��V��鱻벳9YP� s�>��J��<v��7zէ�����l;�-fE7�/�_���Ѭ�D%��x�{Sa�5뽗�5�y�6���&j���ŝS�ߧ�nnă�P|'c|��_�������Z8�vT��j�Ԇ H�O�ӷ7$,���-rO$��G�?n���_T�X��4��U���K����}/��kn��"!o?"�c�~*a!���r�����X�W=N����/Yk���v����M������S�d�=h�c���n��
�4k����?h Ⱦ4u7���#��eO?,�*vۢ&p�
�rl��������u&]�$ɟD��>	۾��gC�a�N�(I�M�v��淵�~����TPSh�kT���	���*[���4��6��j���<-F��E8b|�C��{������ֻ�a��\b�.�L.���]�h�H��Mc7�s���|�o��>�$����ge��#G[_�T^��:��A���7X̨1��� =��c�(��?|E���l����Sٯ�%���8�\Ծ��[�M�&��CD�Y�B���OM��8��/{�^To3�]`�5�[
����t ���3q�G��
<��e}4w���Rn���dx�`k��}���j�A�����R���=�s��Q:���eZe�w��!�/ivc��(6DPG*3T�]��cz?�O�J��'JX��[CN�?�Pn�$�\�B���f��h�,�Ea�?Φ����<�TW��.~t�ys;�X�����9�;Ϸ{F��;�@ɞ�-K�C���l�`��7!= �ŤIT۩��O�����Wq��B|��m���T��l9�t�������4���������^=;)�;�WOj�/H�F��Н�pĕ}�ݿ��5:��e�W}1���3�#hZQ{ ���������`�����B�����gf^�P�v6����{g�������˚��w��p��9P,-��h�R���%��b�!�vk~&^C���vru?}�Xo���r�1# @�?����`�k�����2t�:��������`�w��i�o�>-ɽ�d�=����bno����$@�}!1f�]?�'�X��<F��� *��T��6�ȣ�{5n&�Gؐ�f�Z��hƯ.0���ڢ�U�Z���g4_raiW��q�����S��=��:s��kg�N-�6��t��=FY�F�'��oҼ9&�+fϰv,e-^��uk?���E	ǽ}�xC�`�Fs�U};Y��$��H^'���Q�-��`��PcZ�*��Sʹ����I��x�ѹ�g�{g<rw�����A���څ�c�5c�����[^���Y��߬�=��KQ_�~�����xY}tvC�?� ��ч�:U�x�܇J�@���ŋ���'���Z��f�<�2��˖L�;±�V�V8=w;e��;�-V���l�P.�:m�baW�Թ��l�A瑲�]ӿ��?��E4�~6<�#����6�y��#�7Ljo��ե}*����ľ���X�y�a���S����'7�A�@I)��Q4�'�݊�_�z�|�B`H9|����c�P��i.���e���c6��=%�+��O�����N/�m��{����r�a�!�b�5��IaH��yΫL�?�,xY�~=NUPeT�ۅD����)�g�'� I.I�N��#�f�Ho{�B�xVn8�p��o����џ��b5Y8������i�����" K/��!{S��l�N(�S�m:��C��Z\<�����?�3�"x�q��k~]����񭊗/|�t&}AޙfQ����Z�Ҵ�?����|��k���(��9�og�):�ܙg/��lA�8�4��C��A������m��4Uؾ���P>���/�Bx<�29��ö���{��x��?E_���=d��<��M���58 �s4�A�8ݺVJ�俢��H�'ִ�)����G�.�;��S�{@�e�.J���!�s�؀��o	�q�+bQb��'[�q�h/�2O��;���r��s��/�%~S!i��T�G��}�N����޿��#���w{�/��Y��\�^<;o�H	A�F9�_/����:��>Y↚|묾��b�r�琅U��d�[�Eq��QVmK? ͓�.� 	�����&��{���+���PiN�dVX�^���Y*d~ӫ�Z��]�� !Z��\��xo�a״O��<�I�K�|��~$⸷�'�����R�>M>)��c�:J��V�бs��E���4va6T�K�5� 2��V���I ����z˅q$W�7�����^z��5x���� p�(+�rr�$q9]��OÊ�t��Qtk�%U���|/.<��
c�����aHqޑ�>�T؀�;���]��Jg_���^Nn�Zt� ����O��q�܇���bC�ZF� 
B0��o��^R���(����GU� Wɵ>J�lk��T�X�q
��'{���3k�u/��#���#�?�@�Lɵna��w�����0V.�����(��f"?.�� *1bE�n�-��C'vT9�Ώ���d�zA��Ɩ&�� �le��/g9�vcO�!���C���T�F�7_����V䚾K>F�T�$;Om���r�����}�,��>}����°�^ܱWP����`f�.2��X�;=��vy�Hd���;�h���cr\\����N#���΢;��J!��Vg��tYu{Ci�Kk�#�L�������̇5�v���ZgƀPɢ(��m��6u�B��J~��}o�@�^R? ��.��s�)�dW�3���/~�
�_�=c(�l�|2��C���e1�2������k&�*��=��JC7�Lin�ɫ�*�������{S����;rT~s��`m�MD
�� 6!�ޤW�����0�oM�@����ԛ�A	G\���N�ZMH� nyF��ڦ���PI�����+�ƹQMDhЇ��0���V����נ��%㓯1�hckҹ���̸9����>����G��?b�͇��0����}�Kl<m�1"�3�8C�d��ݍf���x�n���u���u�g"U���F�5QR��� 34�Isr~aw�^��#�Rp�xa�u���\;z�瑧^;4���͌;��s�ܕ:a�	r�-�*��S�iv�|g��z���+��5�r��Vr��HE.��I��f����e��
�Swr&YL��'�;�N;���R��F*�2ӔU$W�+�{�x�tXgK|��Lx$���;o�T�1������'�l�´F�!��FKr�I��$N�B�ڂh��v^mO�Sٽ$�{H� 3va�\fׯ�0���{�r}מ����C[�����.�hN֫!�o�;b&ݗP[� �L�M=h���!U`��O�Ñ����.km"����+W@�EOs�od����v'WI@��/_H�KIlU���S΢lf����,ބ���,jw�C���%t�iI}�(�~$d��b%��Y��N-��l�{H=$���dѠ6��ܐ���=d����[{`��~�c�k#ya��|����n�F'8����Mc�Rs���k ���Go�v�~�=�^M���Z���V@9���r�@�+s�A���s�W%o�_�W��7�s1jrv�$�1�<��2j9�_�0k�j�X�A]g�V7tE�ᬉ�.�\|��r�{:��e�����>�*QC���D륂��C.t�_���s� f��f4���@��SnM#�[��f@�/�jJz=vȆ���-ߢw�m<j�[i�7U���}a�z���`or>Z���f�Sa׃��'�W�CJK�`�f��=bʼ�/�sHN+�\��캤�j���n��܃@İL����� �ىg��ܳ¢�#t#���j���JP��u}�����y�s���&��4%T��lU*Q�!-)�k�b���v�Y��-�y�1�AOq���+^ h���qq�Z9/��*19ʛ��ߓ�P�o!��G{YDr�%�~W�R���f�wT<���k��,��� w��6�L(D�U����r��y�ʶ;��Ԍ�� ۮ��H�+Yí�1�Z*����G*��`�������/��	��e0�ŝt�}�}+]kb �)K�O-�U�t�=JhwO�M�>�+ގ>*�m߃����m��G8S�PPްbȿS�P�Þ���p�`]W�(
��W(&��A����|v���,������(xTwJ	g�4���[U
Y����ϻ�K���tl~I����dx���z���ן���ݤL�o�r-x�_��+�4�͜!7�*����|/�;��~D����m�����KnZqS�6��(�6�f�U&%�vB>S2��y�%����bEng�T�]/����o]��p�
K��v�*IP��*)Zk
�4lh|�8?>ݵ�]=5�KN��$7�n[��N�?�	�!���R�a _˃���  U葇ژ�ܨ�����ղ{�qj��>Bsyf��K�:(!�`�6����D������<��*x7Oh�;S9\��
��������'0�f�L�@�sۏ�_�o��~�|ҴK�0�m�X��q�&�R�G�P��x[�N�۷� u���=L�m elш��7�%O����[,�)����]�����O2�C����ܾD��Fn�� �q[!	wؤ���6XN��24�B�bsd��yU�.~rc��������O�,��f����{?Cy'���p��"}��,K�)	��A�r�e�J�;�E��Ѭ��^Uz��}����_J��,]��z���]�Fıv�an}K����GU�l�|�/��,��l�2٥���5w��%6�?&DO����J�O:�'yO�gq7��Թ����8羿�m�[�~g[�	��HήfY�c>x�����c���'�<�!�<Y���������Hf(i��8���A#�bO�#7��`��4D���9��֫m۵���k�YFJ��.��0�>ۺYs4�;}�<[d��=��� ����4ط�;o%Z/������s������k�G�G�~:|1sr��xk=�WQ��7���u�}�1��N	O���wk�u*i�S�aj�i�;,����[lD�u��H��L��g����*~����o��a� �%Mn��2����~�z�	L�7���m-�j����p��_��lU�!���b=�&w'��QK�\"1�9��Z9���C�"�O�;"\�5����,GMa���}@�K�Z�9qY�X���Or�\�%��^���.���ُ5J��*�ӽZ�(He8�g���p?�1b�6�Zӝ9��dkj^`1�ӓ;,��#$y�֕T5̼]�S��w�����U�̢��z���it�4ZU���ox���r�`���2���A�(����R௎��ޤ�:��:�X���b!� ��[�1��G�����w���	ڒ�Kd�&�0"���X��-B+s2��3:�+�_AH�"x��'��p�82,�*�Ʌoq%��/ 8������\�>ۢ�z�MM+4����{���;<�Z^y���q��Ma��-��D����?�dZ�����gN>K������K��0!<�٧_jZ�8w�T牗�_��)��)ůW��N��J3���"H��\C�%O����Z{G���j�^���9Ztgo��Y0�����D�H�a��Q���`���3�L�Z�O�D9Ml����C�t���S���\��L��o��2 �gK������+]W�8���%���}O� � �X��,P��|��]O�#n��L/v|��Y*��dJ��o<��GT�K=�Vg�5f�"ΣH�D"��:���c��s�	��%հ#)*�z��}/iܵ�Զ���Yʺ����M&�6仿����waͬoS\��!!�P-~r�憠l�Y�"�9����];����ч�KM��|/�G������yji�jֻC�+�n0�mҙU�;��K���7] �DRH	���E��� �ͰIC3����^0�mm?S��5돽$�g�w�I�Ķ�ю�,���_�rb;�i�B[����>Dz�/K�[>�C��_}�,i(��?'},���r�kg{������o��:�����U�O�	{���LA���j�ko����P��m�{g��͇���g�n��,�$c�r�	۴��N/(i�rR�$�۝vX�&<�J�W�Py�qX���'S�Tֿ_j��Y��)u3�][2�>v��A���2E?�F4��h����{/sSEA�����ض$��I��PoK���̣�A�-�*����I>�x��M�se.\+fό%z�Ui��
�5�{�����7٪�ƛ����?�rF��#n.8��k�i�¦�\�,m��v¯��u���vņ��d� ���r�i���Z,7�v�P��?YGW�\r�-�f�M��o�I.��'Nڒ�V}�ⷵ�gQ�o}�g_��^�cWW󉯴�����+�7�p�Ǝ�K>�u�
�K8<��[�d�K�Zy]�aK��� %sv��0�.����㾴#e�H��]�S/��6\θ��~���d���$���Jp۹^�/j*��8e�����JC�"Bs/�۶f����I�����:�0S�F�M�����o���9������ʎ��~��}7�D@#�lI �I�S���M2��������[M\6��)|h5���р��S���N�_�?9a6A��׺Qh%c�Ο�"�x�^7[��q;|��pӼ7%�VV\O��p��㦋v҅��U3�T1�Fd��B�4^R��2j'�Ig��u�#�r)�Ƚ���m�*�x�)\����m{��U_n)�ע�������P�A>�����+��ø�fZ�ޗf+^;"
�(@F��ߣ�M����(�����Z�&2�	���A�1E��B+ۑ�lI1�����E|�y[>%rfI^�9�W	����~n�d%FfI�ig�ބ���QT��a"[�~Ġ��l	��j3��%�昗���{zl��>'?,o�)���Āi�g�p�o���J�H��?ސ�:�z��vruI9O���#$k�9P ��e�H7`;Ÿ�a'��ݻ"+=�r�_��Z�/��R5T�%��Sm[�5�^b�j̟��Zb46��vsa
���~C��f�m��&|P�r6�ޓn/��[�/Ў�G�9v2�s����������z.�ԍ_�&RR���j8'��n�\ �F�"\�L�1���go͌����ڝl�ޛf[7:��#��{����M�y�jcVV[��=g�m&�nH������wwUsk�hW�r,*�6������96�U���DgDtR{�1����4`C���Z<Jw�2��-��Z�6V��q4@8�\��lCFD��g)
��W��	�����4g�����I�B.}_��&�LxƱ!v�wP���u6C�mo	��R��D�llo@�Η�cq�Vn��s��ث1r̍q|?LZ5BS0-WC�<N��]�j�\s�5�uR���a�N� ���Jd���o_���uC�_�p��L��Jj�������?�w�n��vT���zd���`!���<娥K(��P�ǣ	؞�\2��,/��=[�X �v�*U��zX�U��!��E���_v<ңI�r�W{8��a�c�.T5�W�/~�!B;��
�d�����%�l���%�J1)�~��j�p�m,[�y��py���@�g��<پhI�n2v�<u[�,Ko�r�p�4�7� )d�&YHy������c�涾mϕ��;��F����\�p>|[z��"�"$��E�8���&�Y;����^��pa-��ͺ8h.)����irxLSp�-|`�z���6I�8d�lx�[����`�#�����]ƻF��b6�����E@i�==�(kw�L�~�ǝR��;��kI��^�;~�C('4;㞈 9Z��tV���7�d�`@�6�Yѕv<�Kc%�8�S]+�����ʱ���W�o�?��F�bv�5�a粭�%\Y�M;�8b?-n�g���#k�j�v6v�;X�cm�/���]m��S��-��(����V�qI~��O�������p!�L��{ī�;���9�Ҳ�%�e��bܲ[B1δ���͗�SGM�6�̳[3 V�> 'ۘvb�"����褦d�c��T�71,�ǝ�u��-���Z{���V
ԅ9<x)\F'���u�cz�l<���x�+^����#Wy꽮��3�l�r�X�o����ůI����t0����5�CS���j.�-���O$�tR�~���S^��/�XJp��*i�9����f����Xt8e����&�����,*t���-HMSן8��&"x��[�uioM`s�m~�B�Ҹ���pm�ā�,���|��g.=^v���
�����r�wPl��
��7��������:O��]�;:*���X$�C����_�E����$�[����P��D�eg�!)c��gώ��>4��Y狧ݜ��t!�8;��%f5ݽ��wtH�wDT����\/۾�L�a��}�ґ���u�ݚ�T-���PY�;��s�B�k����j�x/�QIn<�̲lI��UM�zU9��7<�����Vm��1�w�����zٸ�n���r�~��(�Z�%���{��G(4Br�y�2bD�Ca�8�Up�8F�&ۑ_�RS��s�`��A� �^�eFn[&��m���]h�γ�]���N3�'iJ�!��爍����ii?�G2�;0
���Qu0�s��`�~��k=���w���%�F�ݤh.i,�����,0�K>�!����a;;>#�70@eM��Gzqϋ���>�pm1)Zk�S�VT���wkr���F 戃��v��11L*&(�[M����j0��-�H��2��fm}q#�!ke��ϷU/f�S���j��U���/���3z͗�������k<!ٝ!3ߣK~�5���l^Dj��%fSo)�vCV��֓��mg�>m6��;���m?����:�DfM�ҁW��c�b ��w�g��wž� z �.����c���|����<��8^b]��苘���D�nb���IV�F��N�$e/@�"7�<��Hl��0a�,�f,��Q5���'_欄:�"�����Yi���`ဖ �J|�	�-�It�|��;��"���.y���跗0�����2�ܐg��r��UO:nސڢ���R��$� Q�$ә�c$A�5X��������n��zivRb)�̔n��J��k�`4t���3ˢ�`(uZ8��f1n�����,�:x�7c�����;�8ۮ��~����<����t�<�u5�B8 ! ��(�A��s�y���	Qd�\7�ϔ�@��Z��SE=�\ך|��-	� �=2B��!)�����:͌����� C�&1�:�v��B�	;��;:����{�De�)Q_0�*�f�~�����k���5>�8h������w�g���u�r%�H*i�=�,��]2W ��%�l��B�A*���]|�
P2�[�@�-���	u���ܐ��ʆ��j[��Q�ng�G���R@p[ ���cɇ�7�A�!XY�D�?���28�u���틙��z�U�R��޴��bhYi^�Փ3��?	��0(���a���P� �)]=�8�<M���|�s��C�� #��7"��~���O�(�?a,{����td�C�A��k�`�7��{����0���b�Wb���H�A�i�>�K��.������o���M/���ˋ����k�D26+�ޏi���FL�O%Ɯ��b�b�>`8��/���b�le����^CMP����vA^ {�,
4�u`���^��
�T�ؙ&Aw�c�C�����vCo�7q@�w�E&�?%) ��I�2>����-!=XDD�1���:d�Ə���G��۱�j���y΄�yb���1Ec�0^;mX~=b� �h����O�UA�.X����b����t�9�AQ�K̴��` ��]9o�s7�d_�nHY��1�M��{HX��󣼛�h�s(�4���r�
�A`9��W���9��^`?6e~r�yY ����6�A�Z٢#D�����:w�]��Pa-�����Y��w���$O��8L��P�9�����p����BY}� ���ΰ� QM;�:1v�
2u_hRK�H�k���/�11��~Ix�Op��?aD,�M�b���ִ[��5�DMе_��s��Q=�]}s���JY�͌�ҍ��y�[��)>�B�|�i��/1�Z��/J���݂7ܛ7��h�֛Cң����1<{�N>u�ӯ�ʢ�P\g�0 V�A��7F?lA+���{�Ý%Sn�W���
��qV�#1{�_�d�pm�� n�fJ��Y��P�Y�
%`E��<L�d�������ӌsZv�'��:�c~n���݆9�W�h"�^�8�é����n�M"'8����?<�T�m�[1�RA����tcQR�؈g������ N�6�K�̯�X�����+����� ̼Fx�03�B��/��[��@��~gv&p���r暣F�������׬��Є�VknH tr�t�I�I'�䲓^:(hk���T/���}aR�I(S�p�~}�@W��}�:_2+܉�U|�72E �]d����%�Gi�0!	
{Q`�Ƌ�)�j8����\b���������� ���E�L�-X�gHl��5��.}|\���+�7���Q]�!�X��	���Oke��2�Ԛ `��d�ه��N�B�!�I������:�K�6?�i��~(�VӣeM��Uk�L�|��(pr�޼M>u���;�/��#3tz����r�%/��0.���O�R�;n6LME��k@Y�n������\���i�Ly3��Tl���H��aߒ�{e}�bBq<��ӎs.�
K�'!��:�-I.0MKkͰ���<d	ͩg�o2��k�Po)2H�Aȶ����ǰ�j��:_g�i���Η~�YI;^9��O��ctk�dcf�7 �4�şx�O9��+@�g���5�1�4����d�}(L���H�R��8���Û��cy{ض�U߭�'`M�w��gbX����/ ��%�e�տ�NW�N���h�:w)�6����;���u�gC��m$Բ�SU���Ι`������Ĥ�&a%��|V�Pj$�wIP�X�f�m�O�����_uE��s�h9�ݖ,�,��v��;��e���pt4�N��e�|
��Jbm/�����/ǿ[��c�������m������L�N��;Cr�#�	�j���γqM�;b6'�q�#t�!ϯ#�=~��yYt�a���\��*!�
8�]-r�9_�x�͘Q�:W�.q;g��L���'�u�8[J�M� �>�`4�䛚Ÿ_\�nw7��;Vx9�x�#��� ۲k��xD3�c�����>dL���?��"f�,A�唂D6�

�I�Hİ��y�����(�a��=ֳw�5Rá��;��9h��-r�� �n��˦�@̦�����K��j,ED�:��h�~�,��x ��P�K�W�/��e�u��Y�t^�Sm���W����|������F��Qr�i�v�����C6��/��#Y\C .�ێ+N
5�'��ztx�s���*-�G�
��=�)�,��tU�]��<~��f+��+f��������E�>Ai3�
��ڻ�,ъ��)~yå$/�d�Ɛ�:�ߘܔjU��&1jWy ��\��p�8�`4����9��v���_D�`���Y��K���SVg�y�,>��H��{�K����0E${���i�H}t ٙ� ��j���E���Oa�>��gX�*�\���B�#�%�lE1T�}�s��Ү���b�+���@$�ye���e����0��dPܨ�px8x�~}�h�O�^��/n�,��M���xx�,�)�����6�U1��{���~�^���p1��[7��=}�������N����~3yP	�����%W��yE�t��nF��.��µ�X��OC>Q#hx �Ϡ%��e|�Q��!�T�����b�R(��El{�i��,�sSʥ�mcL����ȓ󮝗eA����'��C�"9c�:U6"��?�R�'������zx�"u�0ع��n)��G;�88�_�'��/|Ǟ%{f������f$G�0Ini5xZt�m�e��g��Nk,1��W����鳔�I��8�d�
� �@�_@�>P�@�N�#����叽ZjZn��1c��Z_7��m�l���5��,��E���L=&+\�
+�Z[��"?�'\�nچ�}l�4�{6�'�
��sIV�C������y<���V4�%�%�]R�R�`���M�x��ur�β� S}VMЂ:��^=ǯ�U����C��Q���u����򻵢��*�������D)���*��D�	Ҭ����I2%����@S����"\u�h���L���T�Y�#���QBS����'k�Ns+�c)��M%L���W�"y��)~�D�*n����Ϫ_��@7�Z�5囝�_�ߝK�����������a�k�ﮃc�k&�5�-fHZ(��t���h��L��H��-�f��ɠ�½�m��A96��~���FD��c�I]������~�m�lYE�{S�,?@F���T�c���{��ˢf���N��\��6��w>$�jk@P+m+U���W}�(��F��а:@4R6���g�ǵ%Q)J��Z���&��JwT��ؕD�XA�Y�jQS]"�|q�����g>{���@��mu�n7��Y� ��E�������cn�����i�w����C��	�L}u n�S�ۑ8I�G6r�TW���[+@��9{?Il�\\�Kސ�_x���+�0�uJR=�,>��&�<�^E�9	��K�B�-b6&�fΖ��Y�/���5�V�>�Y���3V�[^m]�_��h�vHdG�-�y��k�d.��Ë��r��t�xP
�n������i��.}
^	i��}��:L7�^���@K��(v��'�לڕ05���r\�BS�[0��Ťޱ4�k�Gi<�梈&嘠)ȕN:�^�{�×����O=�|��gB����[�w`f+���6��+Z��o�p�,����ndS��q�6�6S��F:�HtyM��1(�-���S:fs��{�_R^���\��$��VxK����
g�8㎏��Wx��nɒq�7J/q�2W��|���tQ�5�	*���;:����3��������5
8��lX��FB�҃���={ҪM����6ɔTV
@�@�7f�;P|�d1n���~k���X�m�)]��'��΋�_[t�W+b:���aʛv�������8��=%�yy�����l��4�W,�V�"�~6~an/�����y���H$��ᦈb�g�v�G:j��?C�߻w�/Z��*����%ߛ�l�}�BW��ծp`f%�(��@w�O��+[N�������>�k��g�K�;Ae�!�>T'�u׈�L&�J�i�e���a�����!�����ef)���
��(�2)�S�z�ꣽ�+����jM#b5�JzU*%:�q��l��9�����Bn�_2!iPC>^DH�,��lųN���2��{,xm�+��Ǫ�$�HВ�P��PDe���k��K_]�<_VY����ae�Y^�q�;���Rl١��S��%���5<EM�jf�%��|0@	��uP8��	Sa�;�ȶ�欸�%S�p	�Z�]Nx��@k�#Ә�����@��8 �k=�/+��N������xk8��
1���q�Xx�v򉚈���hN�j��#���o�z �>Ь�pz�����[���o�~wJx���M1�#������\W�^��uLg����L��jrF���K~|��u��:�/���լ��9ǴHmE:ӊ��@j�
 ����*����=�ObH5�`�����C��ɧ���Y0E�2�Ol�wy2\�|NAM0}3y@�M�X����.߫�,�9��ve8������#jc���{=j@ݼ���z^� ���B�ߗT�T�7H�m�т������wՎ�#�����{�N�˾|�0e3���ufcOT�Ȅg�!!'Ngeg�;	�B�)n8���i~|x�T��'����Ϻp�g6�~j���F�������T|1��pͮp�r��O�o��r2����Ԇ??,���r�Dj���A�����
��PK&�����i��j�
�$���kGD,>ʷ7g�����5��.��:m��) ��ׂ�?MɈ���AQW�6*n���y���:~�.��yO2`SS�9ց?��Y�J�cBH�ٖw�B���9:=���z�ι2G�ޡפ3@4����qDVy	?J�^J#��4c�&{;N'1��~�����Hto��)"L�=�'-.)_#�<)`ڒ,�ˏ���	fg�vBUL��Vkf$���|�,|��F���'�P��"��f��л��b�6�F�z�@��r���Ô$+frׇ�6{��8���I�c�?1)��#";��ߏR�+�\�t�dDh�!56��&��&�e�J�3��.g0>C��� �lޮ�1F����U$��H ?W��YޝA\��&%���g�ݺk��ԩ�n��k*�)HV���8� ����w��#���X�t´	��<��a���NL��E��4�w�S�cm8䉤��PVD�>�@�V�MP7-��$2�`��&!�Tq�3.�2�������$b�q��%JH	A�K"�gkܿ�6��a��n�} �	^��L�/�Y'�����,�lV@�E5�ݿ�ŏ&�t$�dl�`uR��9�����cX��?�g�T'z(���T�+��Z��r��]{�c	�t��A���5SV˰��ߴ�b��l���k�y|��*����=��7��Zj�M�s&�X��t�!����7^�� �Pё6��W�T���R�/�x6��b��V��S*�ٗ�s�_חD�$�|�K*��ԏ��Jo��N��);Swbgy ��k�Ke��qN��n;Jrs�Z�j�<
&�i;���V1[i�2������U)z�iW��ꋸ3^�:�>.��m���&�z��0�̚. �k���UO��k�O�l���.*�T{��f ��j�q��O�B�&(�����u~����R���l���,���䡝��g|a����{�茆N�<�)�$�$��>V&V�	;�n�t�V�ܧvWU���v❧��9�	_�'e�㉷g ���pDu��N	��k�}y��/�(Hc���Z���Ì����mV�:�}����'�m嬲�"*y���erb���/ �����	x>��L!�g�t:i�0f�s�r����fg���&��h��\=�Y�v��D�:E��?����ĉlQj�@���<7ƥ��E�(=�����H1Ȫ����I�nJ��EO��+�:����|.��9�UvC|�xx^-���8��;<��S�n���<Y���Ǭ4c�����lw�c�}ag �b6*�"NP6���JG$V��`�I^�HL����&%��6}lx��Z�3>�"�j����M�$�A��U�܉vZ�^�i��2ь��̭K�-X�s �/��V^���Z&�J�:�$���+#^�G���f��	$b_YT�v�xШky�Kwg�[�lR��S�C4��!��N�?Ϸ��*�X�d����K�sv��QB~L����&VKu�Mz��Zy��>λ����t� ����|6��k���g��DL���O&&�j�q�I��|Ji:4��m�gz�{��F�Bn
 �/���1m�6Η;�t�<�w�~hL�}e�om����};-s��?�2��;*	q���*���R��'V��*z�be�g:E�����~��ѽ�O��87uyQ�1J���ִ�(n�S䘙t��@;���!�ғ\�\~ %W���
Rq<��������g�k��j���(�S�U�2
����c�!7���m4����ث����8;$�9�^`u�,�xKF�t{��.
��!7�͗��!�yʮ/1]��:xMɈ��T@ՂOA�ܼ�9�ZA����� Гc �	�[L�^�&G�n�JZ����6A�t$��v�E�L�9э�b��Y�H0+8i�;��B��ɮG?40_zU��;�Y�|n��q��w�t�_0zşX��-F�م`@�}er�����������]ժ�U!�fj@����F �d��txO��BM�E����G�ҨC�A4h�L*�lW4'�x6�k4��]�t~�	��P{wQ�������5�Q/E>"0����u�d񸼓'X�B�h�|`�������a�U�j��t㣿Hh��V��� ��q�I���%Ngi['p��a����q�����/�3�G�����o1[�7�(k�m6�� k�tn4,g��i�2����}�SGh�<y��z$�F�/LXn�,bq��7]�R�^:L�]��L�b	�*�&L�D�_L~�;��9�3W�vt��5ܬz�Rӧ3��Cu����_Vmά��녿򉕚��j$��Ӧ�F�Q�"� KY7�Ϫ7����G&'>rs�JrU_�N%}�1��5�[��c�b�ў�m�������ٖcR�dAy�T%�i�I=���<��W�	�l�����Yf�;�I~]�賯��	�HM��� ��~�:�֣��PQ}>%�<��]w�:���h�<���p�;�x�=�"=�l 5�b��>��'1o��82�H[B��ڻ��B�@�5��WV}��^;#I��Ƈ�.�<XZ7��$S,��]u��q�~�ȭB�0�z�Kn'�O�_��*U�	���0O��Q8����\�� �T3���Z��7~`�K�o�}H�<+˃,u��6�XO9�P�ρ�T}��T�A����6S	2�&�C��L{9�3}dnJ�:۝�����;�����Q�� �e�BY阥p̐�A*J�vlG���
�p�q�ȦH�v��=�&2������_�^�u=����y�8���$�̛9z��Ar��;Z�D�J����MLp���f�^A5.��kkܯ�\Ll��o19��1V(����u�EJ�����wP�WE<�O1hNܸn&d�qL���Ѡf��o+���(硴��>�(�_�C8�z'5�Ҙ�K�Du��A=�&R�|�J���I�-���e9i�5�!V���"��s�)��J��Fʧ�U�IF��Lو�`5�c	�I6Α�2GC�w�GO�Ĵ��n�+a��F]�4�W�vwaC�j��6�����z��^�Ifǡ�!C=OhלؽR��T���}��|21�e�Bw{��L�  �6�ٕ׬�� �Rz�{�O��3�c�bd�����z���A�&�#8�~���d04�H��1�7&hx�mǾ�'A��eb�v§h1���X��|Z�j��M�h�=ǋ����9���� ?A�2��#�Qʇ�ç>����J�#�#���)������Φμ2��'`=h0Eu<�Ytf�:_m�O�K�<k�F�кP�y"RJo���	1ͻ����9�==2��r��.���vNc��(6ťʚz�R�V��tpf��vW�y��`���@�a*Y���54X�a*���&c~X�Yy(_���nhy����o.C���P,c��u��4vqj��Uah	^-�˪�~�|�Ga4h5(�-W��U�X��ɝ�4C����F��Ub�)�#�@y���ۊ���F�W95�K���)����a�c������ki�{=faL;�8|P�;�"�d��/�ek�OWj�Ʋ��oy:��Ϣ�7���򢺟ᨹٲBU ���":� }Ğ�}ѿ�Czj��Aˍh�x�ƨ/��=����l;��N3(A�8��Hi3P�s!]���q���n��k�aKM���ӄ\���}��GL�T�U=���U�%�<��;�f�Ĉ���f����;�6�E����4�����ŀS&P�<w�jkPӌʈ��	eh�V�FH�6ֻo���Ѡ+�bҗ��e1�c^=�#C-����Nq/�|jPk9^�L~�H%m�/�0��=9�>�����PC�����]��Fv���O��N�{$Ó�-�졘�C�H9M�@�_�e��#e�A>�1Z�n��n�E�y����j��AD��lA��~��<�5p6�a'�µ��
���v4���S��q[or�rPv0%��y�b��|���e��7����d�#��Og��2�G!MP�ps�tKc2� {�l���	�O���Q;�r܉W�%���&?���?Kߍ2\�n�a\Fk��ba��x4�/�4��P�\�K�D6�#Jn��%��;x�FUt��*y��Ʊz����uFNV�3t��E��	wȇ+傶�}�b$3*ׇ�i��$[!��G�c�(����1��P,��'�hL�*>r��m]Hъ��TUKI#Tu���q�=Aky���=Y��s��h%����>�H�R�M���<�}�zP�9mբ��Q���Gu1w����Ϗ�]�Zu"�	B�^��!��g��c�9>�phr*�������z�!*$�>z,-���Y�4(c47z��xvٸ�X����Zj��:/�������(T�R[�k�J�b5(�:S,�O��E��8fÖ�j�6�vr��#��<���m=�����Aoȼ�!.���I���|U}&�]� 72�|Pqդ*�hI�m���}�mȷ�u#e���H����C�f�w��/4x7y�����p��3�ї�5�3�2*�o�����+\�3)� P���?\H���p�Jd�� �E��Wr����^]��]��o��Q�����֖A��*��rQMM�џ�6Oϵ��W�Q���N���w�)o2;|�I(w��3-p�W�8+���S#Z�O�3�WZކ��^=��`V8ذ��|,���ٽ�&}k��B*̫Mq��;R�r��	L������]p��ג�u*S%~�s��ƻ.��{�l�B`���"�5Q���^T����{O`2��}�(R��_�/G{���Ip�:�k%M�Q{7]�?b��YR�73롔J#�.����L����	&+czX{���P���6ѭ-���6�J��`D�y���~��R��С��C,l����N{�~|����c��s�;,�,p�������헳��y٥�|_c��tz�9��g���(�����W�'7�@�����9����1 �{I�~i*f�Vu(�c��
rȑuf�)�e�4W�%�� c��a�̫�}+�|��=1���3���2�-��Ilb
�O,p�R6�.�}W��J��c@}Llm�l��B���5��5�T+������S��3`����?��hT�e���kl 8T�����0�C}`�jIfj/��Q�y�����λ6��%T*@y�4��2���j�ڰ��K����4Q�jXx�ܱ�k,�j�m��V���7�t��U�2ڛy1�XFH�H�^)؁�<N�H���� s�CfH&�����]+T�3�0�̔��U��}[�����!L� &��4��ֽ�4�A���A��!�g 0��5��L,�_�����9�bb����]t��-�����'s40���:������@^�e~�?�)�^B�<�����^;�(�l(�Ӆ�� $4�b���nW�Ӷ�{��bT$3�OB ���0�3����,?�FO�Q%�ɱ�q�u��&[ׄ����zz�ؖ������I��K��X[+t�8� 8:��#h��s�T���{b�~�"�_��������9,���䇜���
c�o<�@����t�����c���/K��<�+��q�Ql�0���w#m�uy9��1^�2h��۴Ҍ#��^\�|�E�p�t�$���Z����d��ޚK���0�����EKXu�w�?�߄G�;�|�;A��:��z=H��m韣��>l��U(8�~�~*ɮp�I&���r[��������G��*��_����� T^w	�
1��sǮ�J)�����8��^�v���߽=���r?��_�_�?����sP[��*�.׷/ǿ_��!&���-Pڹ��:=F����r���hX�tLp�=z����u������d�R_���3��e9�9�GJ*߹��gY��F����9Xv�ȶ�0R�fS�M�2�Ť�s h����ER^G��t���*�q��VU�Q;���$uQl�2���yό^�Ac�U��W���A�l���bv�Q!� M�r���y�ѱ
"��mT.=���6:˴��
��� �(;C�JP_,+��w/�S嬞B��i�Ȗ-k ��r���r��=�L�1���H�e�~I�O|�E��cF�4�6�6[���i@�$;S���s�@v!�1��&Ű�>�W�+}�9J�)NG繹� bP�|������G�N�I�Ga]�{b�U�4�����ʓ�\�L¿��,�s�k��t�z���qT��}<��$��,��j�m{�@W�p��P�@Vb׆Dޟl@�X#_��U��A����ŋ	G���t\���|Og�R�����F��$��W����%OS���o��R��Sx�v]����?��[]�^�?�j�=���'�X��yS2Ge�B�XD9E��n��A`�BQ�mw��G�bҟ�Ns�6�G!]�w���X����)�m�M�p~OY�챪Y���p>X�\"i:�f���x��+e��d7�)~<D�[d%��Q]I[�98���[������5w�@ؔ*eq�J!�5�=�M�sRW1�<��03�� �_&Џ��.LY ��ňc��}��L�O�۹�YH!��G��7w�������c!+�_}�W�Zn�W��p�n��bG�U����@t����b��_�ۙ��ɴ�/i���L�C��s7���GNt7~�#m�o4^�^W� fC~�����F(���w��e8Z{�m�qX�W���������u�d�gW$�5Q�'��TտR�G�-���\Wo���g3��.�`�����j�bV�]����Ϛ��c^l��Ɣ���o�*���S�s��ş����{n�'�*��Ԙ�/�>�a)ѾΦ^���x���J�H�l�zZݬ��%$RG��&�=�$R�����cg��w��J�W;^)�S�"�.�8?�5��o�]l��%�>h|.:ւz�сMĳ��2��0C?h��7���x;قx-�pYh����a�T�b*P\?"�$hO<�/i�u����2D;���6�7����O��]۸9������Ŗ� P6��z�q�2�ͫ�)��\=V�Eq�z��ͥk���!�ȣ8����~��e�7�~��R7�t�o�����{Z�y�:�D?����o'T���RU��X)!��?�lv�O\l�~);x�+GB;tZJ��e��K�����97:�������-��a����lǡ�8���ˬ~Mb�pԖ_�L�?��,�}4�<�lY�U�Q�o����ʒa���d�NC���7^���֨��_�b9�xc�5�Ju����_k��x)�a2j����x�M#����0F���oP��6��ҷ�ƈ&�r������,��N²i�k6<���G�::�/�\|�*TKz��|�NH�?<���eX.L'�+��bA����)H�oM��T)ᇪ�����e��cg���?ph�i���Q��%U��p���sd%��J���M��s��Y�(�\��a0�l��I���f��V][�x���dP����	�+ڟq�����$�F�Ҧ.D.�ӿ�5���.K�<�����V�\�fԇ�6���!�A�i�2&u����j�Z�Np�/���<��_M.���W��y�~� .Y?��W۷�2�B�v��^i�>l�u�;Qa(�T�f�F�OU��0Xi�V~P��6��t��t�Z~��c�2J�K+Sg�I<mO��D�:�8�+�I�}-�<��E�r�5D4�x�~��r�~�w��z�3I�:4R��ؽ3�sd
��c�I�-��J��؉��%%Vj�L7(g|�ZT|�����:(�L��NW�à�Y;3걩k�4ev3X|S5��0��K���K�r�?�2A�7��W�;y�==��Q�fG#bp����dX�+�}��>����e�f޻�Q��.g�A��S�"��6��x=���v�L�kH�T�֒<u�A1�~��Na��TSa���E���Rn"�2�|���I�
+zF�8=g�����A����^x��g��Ӱ��?8��̷.I�����������w;cL2ǚ#=�!��%Jn��4/�ӟ�z�]���T���U�����ۨ
��l?�1��,B��,a��'m�9��Bb�]�ZjX�3��[J��m�С���D�;��-���8��i���Zq�	7�#1���E��ϥ�o���g%B=+v�+� �{�b��>��B3K��$�R��0�
��m�E�?y�"9�`=�%Y�� �)�t��AѨ�Z��A�P)@�4����8�l�DZ�b��̢gώ�j1�Z���3� r���k�=���(M�wv
�D���ع��Yp6�5f��J^i>���҂MD;-��gB������s�=�;b� ��A���Kvtb��ȝ��{��j���Wa\<�ӻ�Q��]7�F��l�����yVg������3:�CK��������߀��?�}�̔����'�?oI�0���ZYg���D)ѳVd�(�};v<��R�.�uC�IJ��HkqUq��rl~�*�NEW5u~5�!g?~N�?�b�eκ ��KA�$8*l���}�N�F�	��g؅6���
��W��qQ�o%�7*~�,<�e@G��'��v�_3�E{֟��}��<� �.��vA�H7{
�2?�1�5No{V�1/�E�b=�>���y+���3�yl��N�* �F�Sd�A��L��zs�>~�� ����ߋ^���'tF��l�ǐV�y�w�um�g�!��J��L&n�=!�t\���Ŕ�h�{��iv)Ā���O��^�z��@w���Kx�Y�a�fͨ�����۔w/~��ĺ�/JN�+[|��Vd��M��dW�ݙO�N��{*lPR�xY7���E��ݠaz�#h�����I��ڹQ���Fs�����5����7�:���{��6�|�s�۶]4l���1���eyw���EKi����@����G��J���f[�2f&��:cy[!�;�fV>���fޓ�j�*YX�cU�S��_��ǫ�f�v�#~������il��8��oL�����_-[��90@!����j`�vc��t��o�X4��+��y�Y��Kwbx�7y�{�.[�*����K�C��|F��T��k��#t���3�K?e�������Lz\�6#����Ln���-̹,!��	r�bxw�A�r���q�����t�G\����a�lJ�B>u�ϦdN�F� �ƀ��>��ܪY5�<z)�\,����T�����}�!B��[^#�)!-��f�٧�iQ��ި��ĳ$QC�A��g��)�!wA����8��L��V����}o��[M4��� Hv�*A ��r7=�Gct����w!����z��P��؎�ٮ���=�St�֓_j��s���qgl������5�Ss�ZőOf���C�(o'��-�T(�����x��
@����鶍� C�Td	��?�sADx���w�f����&��6�S/�ζ��/��7�v�'�R�IE������_cpn��Ƨ�35������G�~"8׏va�I6�{�sl��CT�ٖ6(�_Ctk��8�5Y#C�<�F����p*L�'��alf�@�^T��}��s�wpJ�����K������D]�672J����h&E���o�������ngy͌������b���,����e1��'��:ej���ᴵ\��$%��_�#*����]]?����gp4�w��k��'�%l��F�������7��Q���2)�����d��/��4���j@3e8����Z�D/v]-U��e�JW*�<��6u�ۙ�a{0cq~'Cf���EɧC�p��1mޗ�N�6��f�����<͖�O�|
�%8����E�*ȗJ5s�m�&ͳd �~ `����]��j�P�(��������*F�y�T��S��_�&9�Ӱ~h<���B�֒���1NV�)��X�/-:E�m�R��uga{Hq)ÂC§ѫ��n�5[��[�9��a���9�c�P`�8A}���$odtrԒ[#ᚾ�G�=�rO��0O�:O	F����e
Wv���l�Zv��c�I�\ٕ��"q�g�a�,A��J���{�
S\��Y����/����ٖ��-[���0*�3���_|
n���Y(���S*]nyy�N3[	��i��!\��*5����>�QVhw}}V}�p"D��(�1� �0����i�9L���G�1~��8�b��%�DV��L��+�{�U�+;
��vv�yd����@U`;�W�a�u9��Rq��]�Pj��
,m�F�j����Ln�S)U)��h2F[�J��!�ԄN�s|nG�)��
f���|���@�c"����!�ޛn:lQ5�3��e�˛h���r^���y�Kȗ�a^'�-\��s�OKZ�`Y�8��]Ѐ��#��ęx�н���i����¤�L¬\%��QDi���7�1zCĔiWt�V�	��z�uR����SK麧�5���B��p���_3�Ǔ���pZ��+��X���D�W����^Q��4�j�Pt�f��V'3��27��L�6i���;nh�XIޣ�K�/͟@�>5���%��U �=r��kO�ݬE�X�Q�<�@E�z�*���<Z��X�J�(z�ō�yЋRu�dԊ9Kl����<�	�Gq#�Q�a�_��
#�ν��T�
�e��D�f�9���o�����r/�������lB����{q��Fc ��*�xN��)���ߠ.�
�Zv����W�R��^j�����Dv���-0I��� ��)�v�r�Sݲ��l9Z��y� �ο6�)/B�I��T�czVa�
f�>H�w�?I���L����¯u<��#Ib�Ѿ
�mQok�ɖ��ȷ�a�,B���ү6ʉ���=)��O4�*�I��A�?�,w�ٮ�U�>>�ͭC�{q�m�L�`� %�|���sB�L�nI��2�v�I:�:^�Q篾�FZ������h��j3M(�Ś/����!��N2|��ی��y��JðYv�#}�8-ĿX;���(�c��I�V�d"���߈̎o���n���3ӑo�t�)��-J�����л��IԩdՅKL��/���6�F�S�_9�U�x�G�_I���)���@[Q�:�J�YȌNA5٤6���@�	]t����8�������B=\P��A�����8�@����h脮�ť.cd*�;���� ��;�4�u�$��v�
�<C=�#G2���V��u�B�����W�O������C*#:���xa_�N�P<)�M���/g{�P�� X����3��Dxf1��.����������T}�ŗ�#}�y4����tY��b�X��e�x� oqS�3U^���J���|��	��	C�4؊7p
l#�?�4!�<�(�aڝ'�S�|�������������?��b��ã5�b+7���>�S�|s���N�<шŷ��^����*�Ul��sor�ƿ��aű\���U��ۮ����WtJC��'�Ej��4�`0�C&�7.�Q�r��A�վ�{�ы�PK    {�X+L$��� �� /   images/aad47697-5cf4-402f-a095-abba84463b41.png�wT�i�6��;�#��*��2c��T	ő�z/�k:"U 0��@�ޤ
��z���K�S���~�)���Y�k\�<�������~��B���_X~��������TTJ��~?wx�����/���T����[����j:QQq|���{�����,�tV�3sF:�R��h�W�VNƆ��|v���dq*�_�����*&a�ۙ3�%>�Or���������~�����~�����~���������~�ȾP��~�����~�����~�����~�����ʾ�?��?|�p~̘�����\���*�Ηsp��"��'�&�m��׳���C�d��;'�G�=�Z�(���/l���d
ʜ������K�Ͻo<�J0����̚��#�s>q@�}�OJY�n������dR5�/�|�(��'�����ȏ�c�X?֏�c�X?��k�'����?����=��$K���8b�+Y���L�ug��J$L�R�(���2R�]�������²��7�btU�謫4�
.=>��~ӹjWS7�����y��|K�]U����Aw<)�~���w���WK����b��yf_1<��i��\b��}`�/.o�U���(��ͬME�������Ͼ ��+8M���R���XP���m��FC�����Ж�D%�w��2K��e��7qoޫǉe�QfH>_'V�%�oכ�)�p{��ڡ`FS��GՕ�ᾰi�)A��+O�`�+�ع����U�&��:��#�S\-9l60�f}u�����P_I�?A��4�O�����#�W;:Hj����Deg٧���S9�C;�IjE"w��)���0	*0�du�K9>�~�\&�A��L�#��|���+�R},����qM���딴��e=W���a���W]zx��K��G���ޑ��:��=,��j*0���{t<H#f"��rT���
t�՚^'��k<�	7��xn��_����8´vsa�r� �߬:ۛd7Wmv��V�#�u/B橉��x�p��&�r��ix���v��Ǹ�#GY\��US����d�8�Gf�`S�����y×3���O
��:
�F��[��{�̱�Q��.Tb.�d��gh���Q��aQ�]��_��|�Ȕ�[�H{�ȱdo�7cγ�5=g:Ԕ�X�e�+�e��ӗ��ĕ������h
y�E�6�G�g���K.s@�'�K��Wk#�\�ʑ�5~�7�/�ݮ���*��Xֶ�1��\����xޤݮ\}3-���\�����x��~޵$��"y���^���=�}M�4�P���=H>�`o��9�/�k��i���#�B#(���z�~⍄��Edt���'as�
A�X�G��ZM;������{�?]�����	��,�N|9жo�ޑӲ�[��n���x.AO�B:�F��C��7�D���;��2+w�}����g��+��fHVotìkP���Â��%��a2�p��M�[��w����#�������!v���,�$�.��� _�����Y��� 0��uW���R�(RN\�M9� �ò�eūع�����7ޫ|w��v"l���ðw����Z���o�yb֏L��ߍ1Tҽ%�O����Z�:�*��\�)2�w����eb�x%��T�O����&γ���hL�l��Ói?�8�S�S�E�C������{p��s���RS������@3��9�j�㉪��5��5�#Q��gGM�\ݘ�v����;��3k�H�>��ZU*z�[�|��>ʾ�Ԏ�N��e{U��`,d�愈���(���P�lA��K�y�
N�#��x6��+��hQ�J���8׆-/���c�=�?4ݯ�2O�1����lP���[^�K��C�h�Wp,�*A��K�d�mx�N��v/�k�cg*��j�_��t�撃�	P��1��Ć��m�d4u��e�1E���?����~%b��m�����P����,�N�N+$�� N0�1�U�8�lX��vq#����`o���nkJ3k���A��T�L�<ذP��#�[��'�g� ��ڢ��$�ԕ�f�iZ�|?L)w�u����2�*�$t]e������"ߑF�!�g!)	l�kʶ)!C�C�jQgm�g�J�'��&�����q(f
v��d�H�^O���f��yL�����HeQ9� fC�Ͽ�]��n�l��̶l�Z�_�Ex�۽���u�)+�
�7��ǵ&jF���"*İ�Q=��"^����°1����g�8M�j��|����g3��>�J(�՜c�T��kt?O�uU�����Z�C��:\v�S=���	."@r���ӂrT�O���3� 2���!��y����3Uحɀ*]Hyd��/�x�����0kBɽ�9�)�\�5�KFM�1).f�V�y�+�[��WnV�9٥_�V��+ڙ�-�o&�gM��{�����!������z��X�Y��ײg2#�T�e&�:;���f�k���uQ�S�
_�j���パ9F�cL�Q��X| a�ev���_T{�+m=>d�_t�?���b�./$݄���S������8���O�F���t#�F������vQb�򕸓���=[�i4��û&���ڽ��,ӽ�!q�}��(F*ka���?dӯTu�5q`vZ���mp#�N��9��-X�*�����0}�������ai��Lr ���mWg���IYm���Z�=mRyϘ�R�4��A�J@ ��^E�Sl���x97��Vƅ��F�������zեh�I	�vt�P�'�%�lk;�~��ɨ���`WԾs����i�^N�ڍq�S^��x�O�)�%���rH��\���l�۾s���^c��OT��z"���}��+*#�K���-�E�p�5�j���5�+�m G�~q�G������k"��s�뙺��&.��-�ʷ���b4�����Gl`9�x,X�#,%������T��Y���<�e�ۓ�WR��Y��V��G]���eȗ��L��̈:��¹�fqoCMa��p�����-l���W� ��	Ѩx}Kn�JL����,����9�k[��z3U	-�w�l,�$	Ի熸 0�Z�	�06�G�i�s��+�S&���6��n��(��@��j�Ż��w��V����6�>q2���O��+��T&�%�n_ߗG���$�$B$%9��H|ЮEP�>�ZF����k��e��}jx`mU~�j�y��/eAf�)T��ؘ��ƻ�,t�������*aBn6��X��n��;�b���ų��u7�K
��Hv��S����T��	�t����⧖��
��,T�܈�ւ_�b�'��k�|���(�i�iO��a�쫊)v�|���ηzV�
�A��h��K�C�wQ�s)���(�+�s�� �2��1��{�f�-�}�I�"��`��]\N�co�W�������`��4A�z�T<�<5�u+�[�m�Wo��.70)Wǐ9w���5wѡ����\�>�6��L?�:'�|�h�PP��d���m٥.�GY�g	K��_��v]	�C�b��`�V����%/��O�灐0��6��O��9��&@��a��� 5��8�+��\�����;u!�p�P����H�i1���x����FZ��ϣr��H�J!:O�����z���`3ğC;<`��ye+�^b�!e�bq��O�t@�*L?�%E�}����|���ia�P��O{>m$�E�D?��ǚK�ӛ����$��Y,D^�K.A���K�[����:b
�B
pAׁR��� ����i�(@��7��z|���:/WG��s����&��CH�~�'M�;Aƍ8�uo���0����"����Y�H��^G�n�fN����#� �ˑf�>���2�c��$�54�����у��b<[$2�{�A�t��:��4a.�k:��p���b�ݖ{[�ࠚ�p�q$AN�fh�j���F.oA�rF�g������ �9�P��>O"��9^�Ɓ��
�%ȩ�#-�M����W'	i�\A�Y��$���΅*�t�"�E�A7�FRC�Lp�Ǚ9�+1�ϧ�����<�o?�Q5�����e/�pm,�oz+�ٳ7܉ÿ9k�E���s���Uɡ�!o�����]w!�(f�cH�����Â��a�x"�i%���PZ�I~��sj�N��7t��Q�X���������'}��ފ=�+@��=k��M1܌��u���Z� �_�=ߍ�*�{vR�v�rMF�)fҿ�,`�m�,�i �(| ����}|q�s���BML�GR7��:/7�^�d��I�:f���g<�,�-���.yC(��qV~�T�&�΢�7A\��Y�
��uQ��t��L/q�|�ZuR��WZ����Q��L�7����#Ō�e뼕�m*����w�2�)
!PU�/W�p�ȸ�B.*��ʆ�6��k������*3�O��B���tx����!�U��z�eє�L�c��)��<���#O|�h(��n���9hâ�ⱒ2s�����O��6]�A|����c-N\/��h��:M&�d�vg��=�f���}5�W��rf�Hg�IW�]�0Iyu�J�[���*����A2�=��,)�v[:{�i*�K���{X'�����n4�n�v����!YS�`�~,��aS���;�"_�M�o�I���8<~n�G��%K�7H_I���KT�v>iwL����r�@����6��J oĥ�|�Jz.14}�1�&�X_������WΘ�|-� `��az�\vޠ�u#MϏ�7?y��h󛼚oREٓ���W���v�>�boxSq�2�?oN앁��o�۰k��Cɬ�I؎�����^ �5WT�M�|��;��G���?�6"�B���J�wt�������#��r����MO;������v�n[�Ȫ�+*�9|�j�e%)mƶ�/|O�q ��>��W��')�z1�_���f����y��B��ч��4ss�\� �30�y�qW7�_��/���{)�.P1��0{����m���M|���y�uMI���zۚ�H�R��$�4Th���O�i�������/{ގ4�] �xw6�ރHʼe�QF�F/Y�ߟ��Hk�ڱ=�|��==���8�S���W����T��p�#ө~���]��aq�|�{|��W��-����!3�Iv���N���o\YlC�Z򹛗��CB�佅�YXގ�X"��ӥ��C~�9
�ט�L6����{g�����JY~*1zԜu�D�t�'Ɛ3ތmF!��$�莶k��N)~�� jM��J�,�l��h>(И7ׁɯ��+!˷̵�%b*ˉ�Y�A-�\z��@OO�F�Nm-�XH��VЈ��3F�O�*����"L��g��c�c^0�5)�u��_�$emo���,G�1�C�q��1�������ݜ�߈�(��M�� x�qlb�_m�&�w�5z�,��C�&�{�6*r�RU�d�ɗ��A�K�C���>"����_���ʯ��C[EY�1�ַ7�vy����(�;e�C;]�Z'
��{�ϛ�W�-6$C2�3�x����93vF�x�OхS��wk�k@8��l(��ǵ"q�c(;��S?L�6m,���0�N]Q���-={ �?l͠�6/gw�4g�+�F�<��μ�K��%%w���TC�n[�|�������ea?��t}=E�-��_z]���kf�\M~h<B0��L�HL*�o�O��0p��.���f��EY�&��������oQJ���,���3d��'7^IA�XoCO�#_Y.�S�q��{tn��2?���p~�0�����w?gػ����Օ]��`��zKd�d��Y��r��#��D�h$��B���=���Kx	kB�)"1�Vy7=g��z
Q��V�=?=�LHh�_r���"����4�B�z��U��"+B�a��o�Y���>��c������ʅ��=��`�P2s0�q��av�z6��m����N	��R��E��a:#n�|9���\����d�'��Y�\u;C-�A��}��4�X�r^3�S�`ʐ���Z�Q<��5>Sb��X�EH�	���~a�DW/�d��-�ŋ�$�ҧ�i9�k)�=Վj;�>麨�1�Д6W �x#r��s5�3u�B��:��w?}���(Kj:�
���U�;~*Q�t����B�����b� �mx�	t���g�m�r��r~8�`��cJJ)7O������V��͇"�3���^f,�>µ��H���O��H�B�Y�1���x�O�0�)�:����(yM�s�.)$�ZC�Ȭ����!��Yܧ�3v���s�7>IA�p+��nJ�`���p��96N*��Q/0�j
�ǐ�fZ1��&��n���W�{�ǲ3���1Z����"�k�!�>C�<�K�Wz�7Nv���«�tbɤ/�")�aw���D�鍊g�,��*�IR��_���Pl����^�w�o*h�x�����A7N|~G/����o�f+݁>�R�d�d�-��d��R�OI�ba"��]&M�o�����OJ�ӡ��[&ꊈ�Sn�ʦ�d�����qrJ�I��K������w�f6�TE�AG��bPH�<<:V.ܺE�hk��cM9���|���~�XS1�C�R�2��^3�}����f�GU��cц|��Y(��+@ 	��4n���r!>���g7��|%8�ش���1����4��TkIg;�c�Xw�3ۄ!k�-��lo���C��0EE���{�!��Q�������cI���񳧗�tVlI�w`?�ƈh/���H�m-qQa�ѵ��wBt��. �v~����������1F��]_��'���E���ψ?�'9���J��,Z[��Y;+N��S�%�����[tE(:8m������g�"�hE%s���z9AO��۵R�֗�/� vW�O�N��P9ϝ���Ϝ�.�Ij��,oT5����bo\v�`�)vk�|�9��-�||_���8������ڊZzyh�G�̀��=�aŨ' CJ����E�N5ȗ�r5��NN��H�.��5rP�r�Bȱ�
�c�R��O��|g9�����BMTH�P>\��p�ˤ�@S���NTO�$�R\ʑ�.��8麆E�e��1�����d�� VyƓz�i2��Iڐ��a�ZJ)��P� �%g�Zݶ��A�gG�w�h.hc��L�~�˒�_������^y�r����)z��U��=~����V#���Az>%���ҷ�(�&��(�������w�Ps�J�c{�G	�5�F�v,���kP�St*�m��rJ'[��Rm��������h��G?�Ÿ��ny��n�H��fr9xG����
���}I��o�*=�F�[ ��L���|z�"��E��d_S��!�|S����'���ә ����k�����A��-�:�Hs5w�IW6sY��H����堯'T�"�"�6�7<��I�zI[Hs�-n5!��+���Ch{{˨��;y��$�.�5w��M�#/��3g�2�[����'�R�y(mSe1���}��x 3^�X'
T��[|�k�Y��IiI��ꊒWO=������6�{c�xE�p(��Y��J-#r[�ɴ�������)�3�.�sװ����؄�ն�N8O����nο��B�� �d@�+at�qeȩm��B�^$�Ԇ�(��Wi;­":ʯ�	��i�(O6l���L���6�w�P��l��V�w���Pf)���D����QΫ*;��#݋~��.-ʹQtvl�,":����{T�� �0��d�k:���o�`L!0��0���D$����ֺ-4�44�jܫ�M0?�{;�yq���}���{,�ջK�c�[��[���]g���OlSG�Dj��Mh����+�����f��
J�?�'d�<o��w���}��3�*�&��j
��g�bsb
봚�q��kO�O|*У&G�J�+����`Gw�j����Ɔ��>�Ҋn�<�����c�ׅ���;-ꗺ�%�!z��`|.9��Վ�bҸ���̟� �3�t�EڕECA柡�1����9!�r�DOM�.���"(�n�JTey8Z
���˩�c6[�ō+e=����FĦ9�����e뱱���ǯ��Y`�Hx��9~��(K҆��`⪥��0�R�N{k�L��wM5���W�Ym������G�Wd�|�o^���M���RXH�%��՝B�����!���w_�mnV'���f�� w��W�ǵ���7���cY��r-�wJf�h�0�c����I*���΅Z*�m�H����'�ls4�Tv��P0,�'ꉢ���`���w�`�0�;i�+_M5��2�2�{�x?���/��|�L�e[n�@8u�.d��'��4���h;����F{��8�%�Ks+1��Q겨�6���O�[��Qo	�l��� �B�+�W�xK�I�u��a�R��7x7�V4ὣ�����/���Sni�cG:|�\K�����W_WK�?R���([�],l�3rMĊ�ڹ�юV�]~�7�@C����?)�`7��}�T���}�,�#$�$Г����N�߳���e��=7��|hx���w����-�"���T���۽�Ǭ�F�a���8�Kz^f���irճ�(��_f���,U[�R�`C�E@C�qY�����ShƸ!�ɸ����_8m�aF�+��a�]�y;�a���?k�H�nh��aޓ:4�	��oIc������� @6�oT�Ӥ
�;��a��p���9F��cu�y1HQ�٧o%C��@q��Zc���3N���,ݥ�Nq�ec� �ym�Lڥ�j	r�A_9Xr���b㸫�0�Y 3I�������rJ�m^J77��m#p�FRB�������3箿�녲���Į���B[x��~ ��P+���-2v�,��@��]�ud;�ٰ���X�i�����k|%_��|�L0�E�jmNv��)x��G-��m_J��t�*�ɻw@~�q7k�4k�iԕ}�l��43#�����aJ�z�צ��~�;RmI.�<9�9 ���pȉ���8���h;K�t�I�z����fRT���U�c/�sM7)�����?���ƹ��N���L�����+��H!�dm�����`��[2 $��U�M�D*2ŝ3)���n�=��xu��pΏo+����2$���eh�z��`�J�ӚL�>#������;�����J����N�S��|��-��'�F��p%�&K���#�3��)ғա]�)�׸�O�z\��F��D�.ϻ.@�QDqe���؇�������؃&��ͣA��k7W����Zqc�����5|��Z�gQ�C�"���������,=Y(���4'��JD2ڹ�{Gpeʕ���.T�x��e��q9���=Ѹ�� ��`It^j�U|����6 ���8����*�`���}���3�R�I�X��/�'�zH�phC[R���0�KPV&Y7�"���ֱˏ�% ���r�'��\��T�^�r�=Ĭ�3�U�P���f�NT�؂����*��6j2L/�P̡!���)��Q4ԒzAT�T�wa������	����MF�k]�D "?��4�E{�a5�e�Ԡ-�ܩ@�R�u���ĄV���A(�^������&}�@���dN��PkY8fVa9������	���'	%��\YUS�Ͼ�eOW.��2��^��B`Dw��t�wA]�{!\�K�}N���J�tN�ƶ9�4�)B8xB�dfo��C��(3�/�}}����'_ٓ&i���|������^&HzL���pB��Cd�D�Y���3����=q�;o�U�������S_ QP�{��:雏YuF�����5u�������NO|Lg?5֪h�V�67�6�p�7vPt\ך��=3�@�. W�%���؂*m�E��Λ�*���P
ʪP���`�
�
�qN�e�פ�<c�#�y4or���Gib�IZ\��[�X�-�Ĳ��,���������o�h8!��l}��)kzZ-��9��khk���O�	PA�\hC��1���3V�>1�����������w�kN��#�Fi��t�S9������/O(�jm��3o�x����=�v��QT|��϶?!m�2��IO~E�	�5ƛ��`�7�w�Y�g��i%2p8�Z��nsp��_<�fhB�VR�=�e�S�[��?�4����5�B�ݎ�'j�{��Z��x� ��'���2ɯ�N�2�g���]Π��`�q>#�Dg�,w�j�r�Hh�o�FG�ǟА�
��s�^��p`�J�:7��,�MT�r�M�e��Mg�~b�Z��}�Ŋ���4�����*e	����ӳ�5%������I�]g~�O���&�nڦ��c$Ռh���/�MX�}���s����U�=K�ܓ׌灋˂Y���c5�m�&RP3�t>�.�6$��Rh�m�c��w��4�d_#��A�	���[c���'z�ճY�f�pׅ��,�GP���Du�DGO�g���:��2�\���0n��_#ra�J-V����.��{��Ql����LAV牓G	I	>|96L�@V	q�;ܪK�m�42���L(xV(��Yr��m��� lQ&"Gʶ;
��?��@)��5�Y��me��lG��~z�{�G�F2U�n��A����Pd�k xkd��(Б��tx���]��~�>�����q���+.<y��fyl`,/��{�a��f~\�]��+j�����KO��͎3{�if�W_��~��/�3X�[{{b;(���<�G�uj��L|&:<Y9$��Iln^a���@,�ns5�����?�'���LG����^��Z-���\ʖ6Gl���N[���sT>���m�C�f��j�3k����x�+!ʷ��Y ���J:��r�0Fذ2�U%���/2i��::�R�=d��C�.s����hX�.����������oΜbH�]�P"�3�OOS�"�8��o#=.;],r��@�!Ƣ�H�UH�����Z��B�4���^��:���3X!�Yx��`��Hi+k=�r��)�dA%�oL,Y���w��@]�zڼ$�2e�1j0�����x�jG"��ڠ�\j�m�av���D�fGG<��_[���Q���Z̐65��¬Hu���2_�[p�T�S�7�3-��I�w�y5�o��y������@�5���y��*ooJ��U�Ie���"A<E�o�F=@]�'��o) �,�㙜p����Q;��t�X!H��ǉ�����\ȫ8��4��=U��<9ꈫ�+a�C��b�Ni�%��#��Ѱ�2�H�k� '~�k-Vu<*��*5`}M	*�8>~/�R�LG�R)�"���u5�͏���F>�����A����!�ȗ��G�0�H�.xH|��Tg�[�6��b�.Z/�uZ:@z~�S�����tE�/����AM"�au<,�wH�~��
#���CǈybQM��!Es�ᶖ0�3����U4��$U�������{��� ��C����M7 ��X,�K�nS�܄+� a��!���ƚ���,60M���w_���_��Y��cz=��~%)nx�Dա�l��n=Dt#o��q#� i�G��-�y	�T���G;����2�U4A��ШW�'�>yr�k��f�NҨ�O���s[M�������m�g��Dq�҄Տ�q��7�_G�ԃD��5d�A5�t���r��`.S�]Ͽ�S>PR�j�u����\���ۦ����5'����d�[KY&m�]GK#hZ!�[�s�g�jX�.�������������b�.{��=�!�> W��1�8�@��R�j�h%YY��2,f�C��C��՝-� D��m8k����t���>�0�;�TL�b���s��Փ-�7�&����r4+�y!3B{��M��%�駠}�ųGw��".��f[6/q�3!v�DW�+�����m�.�UA�?􎅽�dn����V|��)#�J0`&|���A��]ɚ��ظ�廳X��&E�%:�������	��ꏧniIp�D4���}]/�~}�5�3���,�ƾ�د�V���h5�,�Y�۫�f�^�,g���g�	z4'kT&�/]8~���u��O�k_
,���S1+���O�{����yC��8�xt��T��xV�	��5d�f+� �1�F�W���pD��q�N� ����́)��+�i/`�B����E�:����D���[j5����g��3@r�'��o��I�t57�.�ÎDeFY���uG/�zrC@{�da+x��=Լ��E:��/�X��w�Yɑe~x��K�b�ʥ�����*���ɣ~m���88��7�Y#��P�0��BF��^��8�~������M\lP%��W�@-<G|���̾���jw�E�w���+��Y��_�{�{q���ˎ��l{?��=Vj��2������-���z�]���%��n�����z�JJ���ᜎ�����D���gB�Om�f��s-��]=-����K�Y��h���Or��Ǝ�Z,2fJ�O�]�����Xbи�d�׎6���J�,{���}ח�Ŀ<M�8̘,V\��,�݀�ߞMY�\-�ag�'�{%ӳV��5���rbQU��j���i��MX�o��F�M�!��\m4I%����#c��H���z+����k�C�Pvi��~@�N,[	.9�U�1A��Bw��f���|M4*��3nc3��>��3����Ab���Ӡ�[F�t�������E��B�@tq�Sj��8x��DRDBD9����x�\�!��� �W��m�g�¨�~ٙ��:UH�~�n�|���$�>�U]� 8Ưd�l��)�Oו�JE��⪌��������C� ,�hD18ΐ��j�"����c���`v��J����ma˚�]R�������P>~�q{?/�7���r��vi���-�����&;[ړ�L���{��cu���ǌC�`p'a?�����g�������;�Ͽ��Re髷l�4Nو�X��,-����jl��=��0l����D�(7^��w6�I����{�%z��J�*�V��OɈ�/�wrX�^VƮ=��o�^ך/�L�r�S��B)���)*y��W�q$�l/�}&{�[@����z�%V��U#�6�hm�簅W [u�c�G��\N��_r���kz��2<dw�*�e'�q�%k�/9�b���������`���Ÿj�ib����m�����rS���'Pg �˨���xr9�u�v3_W���� ��bA�K��2>v9�H��5c���?�QG�ԫ����v�#�F)�kV󭔸>���M*��*�z��.���>G�t_�*ky�u���H�T��<�1GB^��H�y���}��Q����[v5׉;�`%x�ؙ<m���v3'�7Y�����_�e�m{��6(]�fJP�捊�iR:*�t��g�s�g{N@����5���&)K|a�'�M��HE���d�}�Ez��\��1����c��j�]S��!������>�1f@�%%����z��;��`zz�z�lQcM̛^�w\��D���~�l�8�o%�@0�n�Y_�6n>��mhD�t�z�.l�$ �`(.{%��)U�t)mF2��o���Ãs_���Y�Ð��Yw��3J䪂���ցd���Wm����׏��\�#Ս�h������s9��ݮ����ݴ�,�4�P_�C����m����!{�	��z@��:�+%�K1�RL�3T<�䷞��y'��u�p�8Ǉ&�^��O�O��xiu�1~h8f[�����3H��c �M�W��K?.���Zj��D���L�z��gd��q���y�h�j�qJÀTe!�|�����i�
Rf�N�t
1nPS���nfꀷ�r�8�G����h'���e�)}6�W$j}	��[ �Ç5wP��8���㜕<�w�詠k��,���7�=��y�����*
����l��c�� /�
�M96U�k.b��`�dQ=���)V�5�gUl<��^�F���=Za)�n�+)͔�h?F��<T�2 �!Fo@rw���4
�3��C�`��ƨ�?ap�zΜ�k�jljѳL�yx���v�Pf�����N�H� ��/֥i�������ԏAId5~�$���2j����C,b���;��>�?�����q2�������<�pqo
�X���Ɋ�#��*P��6�S�, W5u�(Ιl3�=��5�wc
w��L��V'���QQ)��hK>��֮ >�w��Mwn�
�3@�����q��q�*]9������4�k�{�O-�y/�G�+:�Y�ZD(=�a��i�'pmk�P���bB�6k�J\Bt��k�oGx�^=6!�G`dEĜ�E���-������\H��������8�N���h%���N��t��"�>�9�Ɖ9Ip��zp#f������3��n��&¯�P�!��$P�����x?�����ޠ�5���Π����������?�u�לc6f e*����儇_v��ٸP�YK˕���GgRW�w5l�>��·�M|��l��(М��e%yO����]\BY.�]�z���7Sc��ٓ'�f�:}�jw׮_�J���-om#5i�*Ė�N�>L��t��>D�9jY�R���bjzM��㷵'���=����L���g��V��H%����O�:Х��>�F/����Pk�f�
�^=!�)�w���Q/7w]_Ջ��}_�tD~o�6��e�bSb�OSNo��O����zj����Ē�e��M|��j'ܓ��5�E="�T5ʞ������=�Jr�Y�;����[���I��9���C �mi�T>�Si�y}�/�R& g�Z-}%[~F����m~�b��|B˷m+��4�*�\�q��+O2DA���ة&h0u6NR�{��+,��s�=�/J�[�t�F����=�ua�9`�l!Ro��y����݈X��f�5x���{p����&��RlA��F�c�#�\��
�|<Zʥ�}��ҹXn����7���_7Ou�a�6#al�d^��(���8/���ҵ	�5�Έ��8���5�L��;̦�Q����o���V����1JzL�zx�&0�ť�6�aa���C�#��<\��jG���^)h��}>*�����
��m���R����'(��g���2R�Zm��t��[��ֿ��Al����o�m��5�Ey���]��MC���� 5��G��u��N�����-Zݭ�v,�sA@ y��	��0I^O��g�vx�O{��p�s�pjM���A�
��1�G���ذ�_ٴl�C]�{qGF�(ag�
����8yt�|�'��[<$h��>����&}�sF�6��]����F9 ���7"�[j�w���U�E�_<�W��
K62�lɣ�@�w,�z[97 �������?i^�hBHKL��BD��N�s]�]�;�wR{��8+F�@h)M�-�\��4�-��v%�Z�Ҩ'zid�o_�83?D5���&����n����N�%Q�e��۔��@H+�C9ȫ
|���͒�U��Z)�3΃1�'>�f9�Wtf�Tz	$m�q��LZ�C<NF	g���h�&�sR�z<�$�s�4-�)���:Z�u����}�`����曒ݯH�k������Djl/���yos`Llw��#��R�Kѵ�Ո>�'�q��s` &�o����r�i�0@��*���s.
2_�%��n��O֭VVR�F�!Iy@�"�m�kjV,6S�G���P��j'R�� ht��U���ΞϏ��sn�H*%����A?zt��l �ރ�kv$%)���@H���LW.~�YV��iп� �5e	���8�>#�G�6sdX/����\[n�O_iS��#B���0��̀F~+��̭�|�u���A��/5ã��w�A%|�*�9���O���?�(f�Y��X��v�:Y��_�E��WO�]�������*2���z�`������ snN�M#;��(J<K��pDS�s5��ZW��<	WtJfW&sL�p,���sOree�D�h�}�:2����FE�W�ֹ2z���n�^B�3Z喖=�je��#�	�nΘڠ���UFS��J��ѻw��<-��͝�J$ �MzK��P�x@q��j��|�1�ܬ�'Vy)(^��=z������10�M#�c�i9m���J��-T�>��/t��t�=]����gD��,�򧙮����|��c]�u���@��S�瞵5�]�����Hv`5��j��h�N�2�P�����)+(�o�}5�|�!fP�N�<�q�RR<�G+�8�n)��O�TYQv�4���A�$z}|��xlmE�[�Gf��/4;�l�ύ���N���ʻ*����Iz��:�7U�PUZ��s�œWfT����'�kO��X�t 6�̫��
=��ڝqx���� �2�Q��Ҹ���5ۙ�B��!�m<Wj*4��K�D@����}y\��
U�g�$i��G^Mva�1��t /�u�M�zM\ q��	�_��8L��ʏ�8�����<�{��7[���"����#˩$ �l�q
�����'ʋ,����LP�ʳ]k/�:E4�k�u�|���U��2�Uݨ�Lo8��˥��x �0&�<�P�Rt���mfU4�׳�g|LM~�I�*9h�� �fA"%@�����>����,>�ZP}�܍ O�톽���
�ɞ��w*�1.���8��W�׊���-� �����t��C}ׇ_Q!�O��+6ˎ���̀78�}�%�:{d�r��jRb�G 2�,�mR*tlxY��2�Dk�+����潂y3o~4����Ti5PLC��X%��x���HpL���K͖ ֊c�u��U8�[t�"p�z�֒��<�
��[��#%7��͎�����P���}=os<c���p;f�f�wN%~���c;���N9�̬I^�(�X�d�[��Zm����$5a=�����G��偁k��h�F��s���j+R���!���1�ׇ���3�T�ż�F�Y�Z��^�+@_S! p���H\u8��bN�Vb:f�T��jc���#��_�(�3� m<K�|?߸�pf�%��G���ʖm_U	�^=b�̭�]2�R�f^�����nD�]g�{ZTBl�ԏ�=���M�d�`o��(/��v��d����!�-�݂،0�����������2]Bu1.&Ք�ǖj+���=�^�OO�6�}�^�{X3��"3��s1\O@9�H����k�� =��L��d�[V��U-4e��.��{"a�U�!�RJ�PS�iT�G�K}L�$�dn�l��YE�/�A�-�Ԡ�ط�L��\����1�e�}$��'SK���'S�yjc������|�zm���S%w�D
��5k�̀#���ɠ�7�n�O��
UǳL=to9�*v�&��g|:�027��[��g;��/�_S/لz��m��b���4���_�)�@�M�V�����RL���I��!�=��	t�x�/�_��P���nM� q��y<�P�wW(60��mKm�k�0�sã�kFT>���.W��cSY���=EQ� x�I�r����e���R���5?��q`l��ȵ�n����q�JuX��T�S�w<"��τ�Z�~ex琊jO/��,"ȒLg`���6��@c�` �/'���t�ݹڶ?բQ�ë��P�ށT������T�]YY�ܥ�$١��E(���:�cӝQY���C�������{�c��^�����~V������z]
�7��K�k���@��.���H��۴�C��":ǎ����Q!�����jҬw�~��s ��ot�.�:�.��[j��7\��܎�p7L�����:�? 'R�x/R����Rݕ���[�>�1����C�
)�;L�R^���+�����=�I��lzw����s���-��2��K9�8Vվs�hT����z�����>�
�2u02�;��w�|�k/�����2o����#�/c�G�L�6�h�:�D���'1 ����%���)/��<_ � ��0�>._�Ɲz�O�F�\�^�1.(�fV�Ր��V�pؼ��lg7�b�O�'vY���ޫ���}H^_�aMу�K;s_{A~=�}������?�3�wK�(�h\R��	&�1&��=��g�]}P���]PVy�f�����E9���4�S�O%����٩e�_�&��̫ϵ(�0���*��?=�u��e���E>�$~+E��oA���yB �u�?

����go7�v�N���	Q��,�r}1 rt�y������ �;
9�%:��8�15�=�>�$��"��~Wp��}�ܝ���W�	g�	@���x�����S�.�w�z?Z���{�E�5��`���u�d��F�r�I��av|�^�y !� L��cL��]y��RV�b��h�o��Y�=&����2����MB+MC6ǟ�z�MxI:̴߿�v��`��{�<ψ���?���0��
��6[���?���)س#���9ɼ\W���pPoղ���o����&>P���qQ�D���n��z�3��-I��c�2/�ʞ���%���?k�ﵫ�[�W��×��nC�wfe�I����N_��,Q��QbY#6�"����s�Y���t`#���*�N�-�����(�`\":� ���-����g��@�I����Xd��mA>ݛ�C�� &`a�N��"�La0�k�JR�"e@3�z���8��������{ۥ����U����Y$���ֿV�e%y����M��`��s��c��M����bΝ�1c�8OӨ!�o��=�t9�+���o{� �rg���Qw�����c�
<��lvǝ�3��ƀ��_<z����F���9]�B�7��_݌7��Y�lɀ��}#F6uB^�p�ޡ��k,��M���c��CW�v��=���Eʖ���u\���з1���Ą�e�pb�Z�	Xjc�;,
n��Pޥ���VǅәvQ�yݢ0<Z�M�U�@/��v,��7B�a�d�F@r��{��Z�2��f���?H���I-����YxW��5�*r�⸉����Z��Ԥ����=@�����>L���i�U�8�s���j�FW�&}�]����� �I?�
&��'#o0���u��!�K&8����)�y
��~a+D1��c�ɕ&L�o�I�4�Y��?�uI2���pպ�������)���gg �����6�8=`A��%���j���8����Q��r��m*X��WS�6ʊ־��2�E�4��!�{���怟�#s�k�K�JRNJ�>��`o��|�w(�&�+�?ʓ�gTN~r�KP[
-W��6�rfT�g��"q�z�*/�k�'BW� �����5bfT������#�ɪ�Bo<�6Ad��%�fv��vl׮��P�$t�����냤���Ñ�N xs��D��^ό4�=܍$��m���m���mN7"\}9B������6�F���^�2Ň)��=�3�J�qs��L�ՈW�,�I	��rK����k�����Sr�6~��ki�K�aj�)� )�O���\�L��|�ps"�����n�����ZX���f
;��7HW^sx�;zb�i�+&=��3�=4%�����e3ҦO�۷�<w>2a�"z\��{P(��f�S�H��YԄ@�d��Oxt�C��%�I�f�~�JP��VLM���#<���4"/�R�z!}�!'A��)6Q'���s����YJ� ���:�ݫ�A�s��`�-l�#,jc��%��b�G���L�� z|���f-Wb��8�iO0�
S���4�?�R"���/��ʮـi��^-��>��MB�j���gApL$^{��?��ln�;�}���X���4����^��p�h�4f\�L���$Hp�~����騛��(�q�Bmǭ�z��Z���C���P�B�.��{���B����R��%���fO���']n��g�U��4�Z�p�5��N��/w��Up ��z&�U����nCyc(�$��g9W����G�{�������;࢝q6�'�3�n�ìAd�>=H)�:.ۏ}Ks
�N���qK�u�+�-�"��۩�_��'���6���6��Ƶ7��4X I�/_9���+��0+���ejql�hsd����l��ݍUwS*�ސOc�i�_��hg��1�~|�E���H�|,k��Ĺ��VBwK����FB<�f���jd���|!�a��-PZA���sa�D��"�SBHN�ﻙǍ��~��8��OcNri�J�A��)��*T �$46�j��U>cu�P_�l7��YQ#���BN@��en���+.�uE�BS�E�E��D��M��k�����ӯ�U\a u�+n��/,d
+8�i|3����\l�w;�{��*��GV%���+�.g�B���b�I�olnpE{�� eʝ�]���W�w����[����!����!�Ғ�'Ѷa�	�4��<+2di�&�7�X��+��{�տw�J����֭!{���E�R�L�����9������z�о��>D�[Z|�X-K�;r�Rϴ����0g�g����6���i`1h['��,�G-�2�e#^�ְ����[���aL^��[h��Z�?i
}�a��Xv��kz��
ĀV�%��#��G���%����.�g�Ɇ|����P���g���}��݀iL}u��m[�`��H�B�z���n��v���� ;S:���C/D�/JX,���2f��)��9~�k�:���.��0^��~�2⡤�T	yI����?�FE��M�r��D����uc���r1#rN5q�B|�C;���|��C��i7Z����c*6v�T��w��wyG�Z6SY��}�#p��s3��`�5i)���Tx�������%_�e������3���r��������c=��!���x��_��2��m���P6����U�K�H���^�r�hk-�d�}D�����bq��þ$F��Jk��75"<����n�)!2����o_���6W.�z�vyV���%(҅��[����-���:��L�V�b()a�$-���up��oE�F[�n�k\\|�{Z����,hi�vd�d 4�N�tݮ�����u�v�x~� �hI;�~�ԣ/=�m^��1V�&qPc[Ϋp�-{zSj5���K��{�}�)��f��Du�L�,��]���n�,���`��;3�GO����`��;5V�����ln'%V��h�_?��&rh�R��:�]�����'Y��v4oR!�vǨA��sBh*�ƞC���\�ʿL���hp�^����)H����U�� ��=�<&M�v�_����8|o�pX,+���҄����,�r�WP��Ev��R���-��0�5|*�{��:�=���`Ux -s�����P�a4�fxز�G�G��4�Qa����9��'���HP��{G4���}�H���^;4��������h�2�i �|�H^�Y��r'{RZ����ɜ���yx>u�VD�
 *YǳomA>A�	R��g����P��x��W-v�[l͋�͕�q|�:�9�?��?�-X�?U��C*�a��T��N�:9��M��f-�q�@��韈�81�m%��
�K�1�7��z�+w�G<�3"J8C3Y��@�U�؇?��Ѓ۔�P��Y�[�&7���Go�yZT��]%�g�?Xw�w�2234)'�ΝU� ��b����gC��o�ϼ��z�k4j�G���ĥ�:�����i�z~ކǺ=8$�,�@�N�����Fj�w��$~l�VG�Vp���*����ej,��^�e5�k����g��8ۯ�."í�	�k"���_`��W�a�l4����d���~�8��ʣ�&f.��>�����
�ވU'�Ӻ�R�r5n4-vhf��G�,�������ЄC��h/r����ݲx)V�X+ɭO��®�T��x�p�@l�����=F*E_w7CEK$�H;`�5���!)�K�U�}j�Ǻ9[���*[��6#��a۫�AJ��h um
��e���]�'I$��O�P���o��3��q���e �
+Wǘs�Q��߼1�L]ݑ9Ԙ�$���+���WC��2c���ͥ�]�.Jk�{���EBR��Q1vL���T5�ӆ�8����g��?�X�����������X���8�6D$��ɒjQi:+
���Y�KO�];��F�����}N�Զ�p�s��x�9Ah�w���w]NU�l\���)�*��?����Z�=������Ig�﫟	[���@su�CF�. 2�2�c�C�&���@���ծ�Tp]t��al�<�?mҘ0���A��]��<@Õ@�,�M�T�:wh���P���
(37{!��M����l�1����u*���T�o�xF�\��\��b�b78���R�Q���c����;K��Z=ɖ��$��e�Ԫ� 姺쭝y������g������!�jO�Zmb���sd�o��-c�q����K����'^��0�sI���G0xÏ?�2.w^��+���:�\�v�g�W-@�<X���,ÃÈ/ˈ;�Fai8��s��1�m�0�E%D_�b��C(@� 4�HK�+�3&4������B�* %٬�:�lJ�?��Q�����p���Ѫs8�ׯ��{����S)�=�]�̮�'�B�+-��?'-@���s����v]�Y��3B<�_�j6�g6�L=8�
d�t
B�Gޔ�S�-a�J�� ͒&vv����I��0.��Vo��]�D�82������!mg�����+�=��ly��T����B:��eKl�,�-+�K�Gc�^}�t(̈́k���M�q[gש�u([�Kv{����8&���s�y��< �(�1� V
���W�N�����g����H�%3� U�"`�g7,5Z�xlV��Ց��ͪB�
ڢ~ێ.{��50�Z�l�ŕ$>��Z8@5�,���&ٓ���sX���$�D��ō�H�C�nva1q�/z��O��y
�[Nu?�W�Es�ΰT�]V��o�_B?�6_�A�1v���J�h���ƿ��Q9R��:8ד�э�h t;��8�l��\����3��vl�Ƿ�	]����;A��D���q��s����dcݽm%ԐZ�gYN��k����#�=����|�ŵ�
���O_����ڟ�\���JI�����Θo�c��w�˕�*�#�}�����Th���r�O��-�@'%6�
&�K��o�pn_�f��:��?9�oc�����<v+8�E` ��^Zz�ȸRh�~�� Ԉ�������v�<� ,�GyG?K7	)�ѻ�O���uȶ��Ӕ�����U�0b���M��L�+�ƁA���kV;�J�g���ߧv�����E���~�&�	�PT��y�����h�з�fhg�C
	�[嵢�B&�g".j�QHo���A�{�ʹH�����
��ۥ� ��������+�UZ������0��,�&�ρ�aL��<�N��f�~�*����Y�M��W�b݅FE@zN��ތC7iNsK$�-֙�0�����jo'Pm��NBj.>������_SC�vP>��R���ǆN���Vj���7%��H�O:yW?��`�|�.����T{V�1�~�b~
��wa�0����9r���g���D��=�"�l�����\�����o��al��_q��fȯ9�F����I����o�PZ9���?wl�e��e(kw��v}��ؼ:gn%��iɨ���a����il��̧�o}�<�<�t_�(��A@������9�K����*/�����b9�<i;��;��'����i}�(l���̩v�և�J8`�Dfc�h�����ꏓn�UlJ��/'?��	�Q9�QU����~��S랠��z�|�-�p_n3�6&��a9S7���l���~����?�`cZ�`��o����>o����\���ѽ�����yCl�
(��ˢrq��}�������;���Zfɼ�]�:�`����²ژ�_��,�@�4�e�����a�uVH"&âfl���RN�{}��q��6���H��E���3>��C�'ݼ�6��cs�W�i��lZ����t�F����0��:8���;i[�;:�oµ�wٮ��3~|���]�ZW�K���!�r�,�	�Bګ�Ġ�^���Gu���V�E,��s����`c�����"���ؾR����r�r���`{H,{�z�����a��q��AۀN���Y��:��$8�&|�~����Nw�͓�gX�g�׮~ϴ_����|�g��R1�Q�	{���w�����e�@T���<���t�]t�����hu�d�8�A�I>'\ @�4s��W4�>��{�iK�ci�G��\���T�W�U9Fߥv��3_6@��~=h`���h��PuX+�����"�4^O�ߕFK�w�"�*)����Ӹ8�����\v��l��k�&�[B�����۹8:L��o@J0R���aƩ�l����83'��6 � ����	��,{&�Z�W��TY3j�.,<p'e�'� k���|���r��'��/M9��pɛ���,���A�&Q.�2����3�hg��j�m�I�V=���t�\��E:�M�%�n]�S�е�.=h�l�<&����\2���j}�p��?4��>���$��>�DVIs��o;{&��]�,kbZ�Ǹ�V�b�{���i�N�]�=�a?Cc�J�k{������֘̐Wj2]?�m��][��t(ЪĻ��E	�uNq�p���D�CY/@H��c����v`L��z���>��y,���+�^�dP�h����	ԓ׭@`�Rd���$��؈K���`�v1?�*�c�����[�{��� ��P)�zx�=]&�*�Ze�	��v8kJ�H��V���Y!��Clܛ���.g�;¨�eTo����,�=G:���XK�!®����s�U2�r�d�-�
f�a����<�3L�C� �Cc��>�бس,-���V�Z�������3	����{�jl:�D���VΫ�(�_
�85őc��r! :��k�I�5h��+;�H J}c���<�������8UhS�
Ģ*�U@D��y'�8s�c_�}�L~էn����Q���ߨ���z���^",�n>�To�B��ͲvJD��ݫ�% �o/�=T?�Ϡy�*:w'��l|3�_�[�g�:rX���`V"��l*���3�X���ۯ@Vk^ĳ��~b��4ھ@Gn��8�]/�6w}"��ԟ�ʩ���'<]Ӎ�l�8l9=��;Fc=�2w j�~u
��,H�B6�����K_ʩ���Xc'=_�@Dxp"Pi���܉��ˎ{��K��b�.�"���������n,�h��o�Eъ�� ��vMi+�1ʟ	���9��~��ȉ�5�I=;�;L���L&�~'���UcMѓ�H͜{w+��E�$���G�t��l����06�a��:�3`�����Ʈ�40������a4_���Z I�(�A6ZƑ��1�/��0�ИƔ��|��_w�n�d1�0I�E��hcS��ׅ|-�ʟYeE/�P�Y�M9��C��3�=���>������e�����x��-�dc��'T��Z��Րx\=��d9"���z�Y�;�R��Q�,GD��^Q9׀i;D�Qt�0�5�F�#����W��Y���W��R8���){\����S�z��K�z�
i�.F0���V�����n��x�I��As)��߫��7[26�?%�6g!���Y�A�D�OL�Fb�Yuy�2 F�
m-s1�����/�;�w��$sX�VOU�q�8�g���>L����ż4�II:L��c}kܻ��I��+S��藿��S�.D����md�lGf��>]0?�Rsl����L�T`a9!?���AװY��x�%j�A
s��:��g'&�'��2�s<�������讎��<@Xeھj��\:A�P^n\ނ�ݘ����D,Ml���{�������z���n�����B���ZB���9"lsh;#]�~��������^Ċ"/R^m_pQ<�C�wȏ�[c��5�[����������DDJ՟�3y���=r�h'PG^nx_��������/BǥA��M��b�t#�� �%}���6�E�����V��n`�'���:��K<����;�E���d�h��<��eX�*Y3��G/���mB��h��`5�U�h�D(p邕(���O}�C��T�jfɊ��ү+�I}���D�C�ޣ�`�j1l��U�	"�� 
�=O�QH��eѫ�`֥$9s�z5��VuE~��%�-n�խ������wȁ%����c�+_qAt��o� �m����"9�v`�<@
����!�hR4��H��qIz����0�g���6��%��?�wf�߄��Ӻ�=� ��� A��ů�I佚�&���˂,��.n�V��`�j,��h��m�����k+΋��%�.�ZJ�
v�x��q]�E&KBB��]S��4���
7�:n��ߣ����;��VSAY!�B/wTx���$[��:1k��Ł�DU���SX,��o�_|�j�/�T�6վ�p<���B��y��c�Y��~����uL|��;YХYy�Xn�T!2Lf����.���K����f�V|�s�A�[�B��L�x�4��t�dX������Z���4�%W����w� �f���<�O�o9Ԏ̟�5e�x@붼�>���=A�e\�h�pV��)`*�0�o�F��b�B���t��8C}v6n����=�?�{6���^��I`��ͪ��tM���",V��c����wY 0u��|+|��ց,�A�y�u����zkͫ=oU��5]//VWQ8�`)V��a[?���8�k&%F}�����!�l���㥎ڽ��7����I����P���Й�Θ�2=��"'g��Jkw,۫]��&CH)Q[�A���m���{��^�����C^���}ݵ��P`Vl��Wn�y�d,��L����������T�0�����_#��Ǟ�,�%`1�pU�T�YRآjO���� h���?(Y�������yc�\��YX4}����/>�^p��j��r����7^~nw���:��; ���V�,�0�@.#��|�ݐ�013X)]PY-ړ��xs�<���ݸ3z>^,hdz\-�o32��Ǖl�*���!<2�������F7�1m�F���]st���F�^�%-)��$�Lԥ��jQ9�I�ݙ{b���6gD�R��设$wӠ�b��X"��}5�g�W�fk-�V�#3�O1����L�ح�xz$Č\�]��b��BK �K��m�0�w�q� � ��O��*&�4\?Z7���y�����<�\8�g�n�w
U��V����r)�r��P[�=�14����
=�h9����G9�4Ϻ�`���r�Q�BQj�_��L�eٔhV9?��{ �0YU�n*��t:Q=�o��g���lDu��L���k�����<�ߒ�7�/���6p?�U��f4���`Ajʼ�X�]����?`d5��g9<�����7���y5�UI�{-��|R,Ψ�8����GJ]6����9�2�I���``�v�ی^ο�6a1{/���&��oB����LG�\͜�k��m'+Jp���v������Y/��c�k�k�'
[�F$��+:��p:4�@l�ޖ	�Լ�tt1`�ް�p?�q�/����f������,�t����Hv�-y��yJ��e7��թ�� �ɓ^�)����E$���]�����Q.�p�Rڷ�y��r�j����� Q8*'⻲s��7T���ZMM�dms��ԥ���$ș���q7(l��w�.�@���׻�`����D�[4xL�h��]L�У��{�F���u�w���H���u�����u��S�붿r
c"��o���$���a��鬱�u���`�˃1��M��f ���G�ۋ��B�"�C�|�+�qs��+k��ͼ܌x߂�w��
�ˤ�N:�(�zx�������iwW?.Z���]T�r�dx4\�����u���mz�]���ٙ����Q�BC�����?K��~��y^;��Z~:b��s��O.��d�ܾ�x��߯��{N�<m�6@2�AH� �=�y=���Oo���Dk,
N̐�:��}d�y�t�`�v�8��M�<�$�,[>����Ҥͭ�FV���$}�'~\�����ӊ�i������X�F����m�tؼ��IÇ����0�҇s_��9�4���q��]U�}J6qte�;�E�`sa��i7�mYp}S ޠH挺R�����I$��G�?>���1��D&��Ct����{W�^��ZF�Xۏ�hh:I�2��T.���tp �;ʸ$;n7��C�.��fֳJ)lBy�P8�\5s�"*'�Z.��_��A$��]��bm[L"Wv�t;�vu���L�������Qb�Ʌ�{�:���^��21��0� ��y#MD�}�e��ٚ� N����l�к?�����T�E���P�]L/8�:4z����l�l�Ʉ����((���͉��I���:5�>%�X�`3�>�.�%i����_O�K-�11���������{�3��Y#*�Ի��\j9�z�fWg�Q�7���U&�[�Y
*Hy-~��so�s��χ!]�2�z�>����I�s2�,��g�qÂl�o��F�>����8�=�aa���q5!��Q�����8���f�?�VA)X�闓}/{V���&�j��{mj��'a�U.N�����2���i�h��WSm؛A��i���J����7FN�@���
&}��w��w䊔#��:W1���=rNc�5�}`�G�f͞eR3�0_��ED�3_���������@D�T��퇫e�Tq���`�{�����A>�v=��k��ށ��Zf�VH8��B>6���ں���/���Q���ݡVy���=�[yS<�D�ZP� <{�-Y�/����d?j1�X��j�k���TL�s@|�m}qq�� ���j�Xg/��PHr�WƷַ�2;�鹖�=`���%r+�-ez�m"P54x*P� �QÏ������U�g�� ��+H�w�]u�B�:4�ٯ�ǟ6n<���5rRR��R7��J�c�XS�%%�'ٸ9�7���,/�)c�f���$$( �l��n]"�=o:úH��`L[>TY���C|���&���OԘ��RZu����"J�n�F�ÿ7�`��CA�<���]a�]\�9tԄ+>�|�`�pfc��	]��A:zǉ$2v8v/��k/l�p�'�D�?�lR|_8�_������P7�o��| ���	�����z���zdaK�DS ��W�u0�H�=wr28g̡�8Xj��+	�nT-4D���8v���E�,"8*X�	�9��}��t~\4d����2��Phrw�V�}#�g��ſ�.�us��f��o>򀿡���\\�&�R��b�����8��%n��kA�F�ZO_���7�FJ�v�h��[O]X��\��3(��O�o���eP��8J�����'�~�*.�{����� �$Q$��[�\?�e�zS�VK�w
��YV��؎��rYc8����Ԃ���?gʢg�|e��4���ER�m1�Ѭ���W{����8 a�.d1L�1�
��I ��3�MF�I8a��6%!<~ӄ*�&��l���ģ�n��U��M��j>��q��d�!��~���O�6�����1f"�oɁ=��ɴ�`Nda{���V��8ũUE~���s�X6ݹ=�4�m�����I�c��&:�
KwuՒKj�=`����j]��n�N�' 3YubyǼߘUm��$��`
Z��ɏ���K�G��,��U�`$�C�6Rk�eH��Q��<7��E�oz�qN���5l���3�6�����ډ�,-)��A��������'e�D���|M � ��a����VSs�A����>�N֖�/���'R6�FO�~��Ǽgy`��U���>��@�g�oz1� �q��a<9�a�v'|����GOXPܝ�Q����@��1�IΜ��c����
���cNڟ��;+	褄�MJn�3Y�2����r~�������+�R��>��`��{�	!��˸~�Z;ڭ]�	����<RZJ~�� .Y�!�=B-+h��x��֎W�J�b�168������n@�4ܨ�����N�3��7g��Dө���O�&��/X������.�
�E���ї�o���?�ү�0| ��l��ݜg@�{� �4/_���Z�0�J*ϳ�/���>�1��r:��[Pk~E���Nɸ��Ԑ�G4J6MU5��WC�\�ω���U~	��2�֟��J^%����ШT�?ljaѠ�w ��N\�E���6۴��OJvl�Cm���iҢ��W��
ɛZ��IRh۶��֟nTn��5�� �1�	b�|�kq����{��w����L�������|�.���_��4������Q�;�
�k>�[n��k�� d�-��>~�^�z�2��gƇ���UH�RR+_�b�ڇ0j�6@Qv�q�-�c�����#���8��[UĆ�
`귂!s�#S`#���[�Rn��_S��+�H��v�#b!w����o׾#�gt�������]����-7s������@��T}�,��bzI�G����ו[z�� s�U�ˇ��P2�5�Vs�hW����e�>8��c*�bci7�sgG�]m2C.��bi�U����ԔP��ɺ��Ŝ�]��+���K��5����9�����I���.�r�/f�1iǣ�i0O�i�+�ce���.z~�c��U��>��wZ!�ܑL�|�w����x8yb`u�r��a��}`D��p�%L�2Њ�ˋ�sj�����(��iñy�б�9��~�u�/� #��%WE2i��j�w�/}��"�*_�p��J�n��
�1�>k!@�v�(���>�a��&�;�wQa;����O�'u��
D��M�i|L�ꤗk��CL���t�& �;�$��� ㈖6W�i/�i��({G�]Z0�����_��v5v7Se{��bu#���r�[�%o��t�~��M�<��9���w�cb��g�W}�ϤYw\��i3�&���=0:����6���}'���bC���l�g��V�\�?�qC�r����S������ݘ=L�]�y�-y}n���_Y:���RQ���
F2����8�8~:g�i��r��A����ǧ,-'�f�Bh��I��=���k��[`�~�|H6��G7cFj� ����c�%dq��#Xc��.�=������_ ���� �zm<�9�n����,�N6����S�Nu���KKzv�J2���Ĝ�{��Ts4:3�),L������O���/�����aj�o2�9"���^������>����H��#�R+��]�i5a�k�b�����Q�Q�݆@mw-h���w��r��ӟ~���U3�0�e��<~_tO�{ C�~�_)�� 3o �R�G5�јN$�?/p /E�Y3-kC~��8���1d�l�xܠ:��_�}̧s ��c5�hIH���;�P8�j���y��Q������9��J3�����P��b����pS��%��Bv�'yo����  u�G��=uP%X�����#��Ƽ<N3JZ]��V#�@Ka7�����'��z\C���0��� M�޷�m��)$��DaϺ# V�';	  |������DJ�JI@��/&��o�j��j�T,��K���xƄ��?���|h���s��ˮ��K����7�T�Q1��P�VqP��+A	���n������V�@�U������If>��J���a���a��x�u~�w}�@�u���ԣ{xg�����t�_\�U�������%r���sTGc]M�7A6�u���c��.ԞcQ$uu���:Cmc�ʼxh���vM�su���p��`E*}3�Ak[hV�_�d�����&u�V����]�ov�?@�3d��W�n� �
(�5�̖�u�F�L�>�u�)�}���@۾�v?(P{?@Lv�)�i���Nw�0�;���$Z��U�ǜG��cO�`�����YK˨�{`�J��������:d���?���xG;�dP�����]�\�������oz-�h�#�{�)�B:ߥ�V�KO^�@g,�t���?�����/A�A�Vjb�'3�����t	��R�1�����c(�9?�.?���Zކ�'�{U�S������^�
�5��l4��U� T�ĺ5l��Q���[�]���2D�nyW<A3��J^��_17rf�O_���@����,�Ժ���D���XۖŦ8v*�hA��(���S��ʾrrէ���j�Ő�=�wqi��G�5����f(n}��ܕ
�t�[�P<xk�e����TY�b��eT��'�X
?_#�}ua�vWG���;0InYhǡ���Q�O#��{%���� �K-�@3���x%�m+�����Ղ�YbY6c�h���Rlً�JΥ�Q#a-W�1Xb����6�@�S:/7@�z��d��Q.;��I/�<������iW�W���e�! 1�j�H ���ᗡ{�'�nU >�ҐHLf-F��2��C
����]��3�Qs�C�c�n ���s�h�nw��*� i��IIYa9Ǜ�����8�}����Qwմ�Y[����N�T�ǔl��^4�os*8j{I�i6y�f�J�2�>c����%�Y!��������~z� ���5W�Z��{�jg�B�M�c\�N��!��qd�@��*�ul�����% �\��9�d�u;LS���4�J�o��L�6X��I��֒�t	K�ޚ����v��pnlO�:���$�}<��X��ٳ����^��#�Vb��W[�v���`fά��ث�8��4�B	��e-�u_�&�a��Nc�V�"��8��w��0�&�����I�;}I��a�J��1}=����]*��p�n����o��i���7)CŠ�U�bM`�� ����#���������q5ѡ:_F��,��z��O� 8{v�WO�qs���W�̆�����k3�>�GG��_��i���j !X<���9��A������d�δHY:J%,nU��cYk#(8殳kI�v. Ps�G,�N40�� �$���|�,B��������P�<-��lC����������?�J��;����}��u�l��%-������w%3�Y~cӆVXMA��e�Nw�zL�n]���{��O�6[�M:�Id*�v����)��Hvq���cz��e�֏�� D�ų�ߡ�+fS��(�
��%]&@]�����,�m�0�;r����+Y��{��ƃ��ONȿn�jo,�d���?��󂩕Udz�"�"r��9LW�$U�A�+�����ٌ�:���ߡ�8q1��:���%�R���=qӐ�0e�k�a4�l���[��솮�Fk(oU(���~�w��;���x��?�Au�Y����%�ٴ��Xzz���#�a:��û|h�"=���e���d���W�°�Լx�0�}LG�$��P.(Z����D�'T{�o�ܣ���܀g*��RP�5�2֗L���;��)�Y���ӊ�8b�RF�}���J0��	��h��[啨�Ͻ�{��Eq��3����h`wd��_���@꬟a�����d_]�$����n�n��ƙ�?M���=�L��|�H�٠WZ����Le��B\�*�m9>�*]q�J:�nl�D1�%C.ۘO���D@�k��\����jA^(U��� z���h����W�eY͜���/�f&߽��޼.^U&Ņ� OQ���T]���Q��2-Yj�Ļ�RW�WVe�&��������V�)t"�U�V��W�|-�FzZ���lV����}�3P��]���<����ס
���ր���&^/�R؋;J4�q��>���1�-tU9��y-͟f��B�
�Tv��V�z�/�K 0b'�������F�ҟl��6f�SA�F�� ����(7���s9��̀'Y坯BY�;^f�'#j����	۩�������*_cƋ��5�[�9jM����6t���-���F��1��`ʞ]I��/@�ٚ*��xKdSu�2=}��s,���_j��2,�:���Z����L�N�Џ�P�^m�mڍ�x�1�/]�4l��̍�zh�=�,�Ad���&�w�ܒu�������Eh��t]���Ը�__��3)g툷�1bU܋��G���0��<$i�ao�� ;��$�ۧeX�~Śf_����?(n/�(t�1BȲ�fu�6}��Tc�=��- N��?վ簯koi��y��HQ�4��a�j�y�c�t�X~�ϕ3��B��Fc�%��%�R�y`(��s6��g�"�Ƣ��VN�%��!D�GMpgک��uv�UQ���߄4JYՉ�'���Q 1�����F�ۀID��??��y�ެ|'��� 7F���V0�Sl,}G�mrb��$�u��>i˂�^Y��6�{����0�8��O(��Yd(9�����N>S��m��!,)��Y���k]�E!������{iC�l��l�2U��+�,L���vv�����S��%�*}ߍ6�s��PL�w�x��IC@��8�tx����sڹ��<��ޖ�����,Z���Le��ܲ�V��S7
�<./9�_K@MSb;Y3�F�F�[d�@��9�Y�ᗁL��&ƨ��͗7C����S�����7<ng�\p͉����ۢ͒��s�`�\^��%&�=ޗT��&�ip(�ߜ��a��%�kw��cҎ�e\�8��l���s��e�Ia7��tJ^������wIEъ��I��Z��~���6neH�B0��嫹6�tޏrrf�[�A�-_M>�M� $b��O��Mr\{8)��3�@��{��ʐA���Ŋ�?t���xz}��6� �|-����m"��NqT�:w})����\��-�c�7���=^�ZS5K9�]�X{����e����$��g�i�u]�Q󳞁�I�>zҧ��vh������qQ$��𸸀Jr Q�]�$Q�� �"� 9���s�AQPI*9�䌒3��"Ir�4�0�a~U=��|�������Uu�9�[��7� ׼���嘪�Pg%�����\��m����n�-�{���/�������"N����S�����,�ŉ��J�D��Q��`�E��@9�Ԑi��A-�$r�O���te��j��dEհ;�&Eu�5ܕ�ӏ4=�G(��(�+�cx���b
��y޿/�5Y������-�ݻ{Ms͑,X���O�p��?Ű���&����T+����s'	��wq�t�Ě�6C��0��N�2i����)�O��p��1��$��JE7g�mѲ����GqVI���Be=(��������-�k3`ť��Ӌ�7'�����*��J��\�K�9*������W:�R��O#]TvJ9��n�+ˀ�D�B���g��K'�nE�<2&U���h�J����DM}jsŃ��m�R(� R���Toh�����^F�s�;A�b3�n_Z@��
�&R��NͩX�tpM%��S��DP�V�zp�k��B����C@�M]~�X\������p����ƙU��ߚ��\T�g+W�x�����#��Ovg?��_�r���?bǕhjy��SE�?�#Ҿ��ʞ����q�������fU<���y?ٹ��#����YO�럊ˬ��!�wh:cgy�V�;�c��:?�R��n�!�e��l�Ad<�0ǃ�<��Q��*�7�jno��
�T�Avd��������>���X��rr�ZN�0��xF��u2���L��{�3�U�5��kBEsobBf�3gC6�s$@�8��&�Y!/���'G���O��WGG `���[x$^����*�����E���E����)�M��Ծ�ۼ3��@g��l����Q��!�:zb�B! ��%��!���tw'Qe�!]j�Z�"��*|��'��:U91mC�zu�e=h���1�<Ms����˟QF��]oDX�R�Cޥ�e�����$2V~���x5j���<#7s�UÚMT��T+���)6���5X�:(H�ฎ��*7���!ۏTn�*�{��p���������D
!oр^�:s�/��a�P.L�j�uX����ޗ��w���_��C�w_�n^��Y��	����%�r��х��@�6l���(�T�,�R�h�y@�}���g�.B���'�ծF���%k������xo<��O-�ziP��:������z��ӝOa�"�^To�*RNqd}烮��nX<`}�O��3k���QJyp���ȇ�S�&z�X���d(����wǚ^�@CD���6t���$nӛ{89�w��acz�:zN�X��s�|� �v�1�,$9�dY��k���0�O���Q-<9��qw�X�R<E�$�h�W6ܮ��|e��ˑ��ٔ�瀼t��J�2GL�-��T�	���ʭ�$�+e�*u5;��R�7��vܕOfwd�������:$l���Kc%h�+�@G��]���1�����cp� K�	��K>>'3?U��YleS���Q7��a��ٵPk�Y��^4�/�B�{Ng����;�����q�MSٱ6b��1u��f��m��Dt���f��;!�x-i���ܽx�}���g�'�6'z�)�_/�4z�	~��2�i���`wP�r��BY;G�v=���3FO��7�D����&�g�R?��j�|_B��@AN�0��xP��Ձ����β�d�$�5�{#Z�n*Q�cԯO��8i���ʍ@n�p��[\��'>l5�ӥM��,
8��b�Sӛ"@cd�^�8���|�H��#�RLfn����5%�^�v�]ﾏ�2���N��[si��^��J�@|�wծ{5�BƨREm-�^A�R,v��_
�GNS�������8��_�v�&��-OM/z��w������o��A��Jޯ��P���G��/�X.dZ����ֶYD1��τ3;	nP.E�d͵���@������v#�=K��e�(���nފ�A�ɹ�z�y[^�H��gs���|�+���z�[ӣ;��d���7��]�I���a[�S�7�R��a��H��'�)�����N��[��tu���.�vegg"����!���O�Z*I�zގs��`p
ܡUv�J6",��κW=�6�c&��p�����Ҫ,첥���m��9�NVҸJ��� r��.Zx��!�����{8x�Wu��PQ��%/`�VV�%��"T��N�'�7ÌR[n�|������~
�{uS)�vU�y��Kp�8�b	[L�vp��A��X/����	9�m��i�Z����\�L��t�����ˡ�"z{O�ijp����.E���(T �,y'���rv@|���a'/�Gߏ8Qc�	{g��n������̎�*/v���Ce����$l(O�~��<�O����x�Su�
V��)�+���������� �JN�ɖ~�6�B��5�G���8�!yC�f��SQ�h(Z�T����-;�j9��7�l{3����*�Ϯ�>�q�ZB^�AQ��l���	L���ލ�ao��H�!oB�Y�t�JhoV����넕��q��ZbHk`H����09���~hz�d����$�>}��k�"�W2�> ��M�2�6L���qǤe��G�6=�y��}{Z1ٵ1��b����Ĳy>���쐓���wqq����f����c,!C��5�.��e-������<�+Y��dl�^z��892��KiE���6@g���Wfm*/X�H;�����
 �3�'�;�C6�������If����Ip�R����fa�ލ�����s�#�
�I��(�Xi�����_�eQ��"���ٍ�Y4�"�{�$�����3t5e���l�ӄ�dB�r��'|>�2܇��tZO����vUR*��I���͛� ���M�uq[$�yQ����k?x̋���bzGdA|�16Eԉ�M��3iQ����� ��_�硛]L����ʙu��B�ԟ[���]�����_�%ZI�U&|p]�b����<ؿ�3t��!�}��-�&��_�lǻ�:�.���RN�+���H��U��$Nu<���n	]M"xo������F��g-�������.�/l`�k9�ްz
��|3�9@�ft��r,"g�����w-�(�\d��|�hz����o������HU��T����[�u�i0��-;��p)�ߦ,������{K:��)^fh;7�>pTLE�a��>cR����>jԙ+�O��5XK�q`&�����9����?�^Y�8t���e���v��Cр������x�\�Ârl��G�H��C7��{�})A�y�Nթ�`S�ޭc���ǧ�V�;�3Ww��g��IH�P��/U���?��pNNn�m��+`:��芋��(�|�qʄ*�TS&$c��l�-6����2�>��vܪ��E|�`ٜ���i�2t�g��=|_CFT��7����F����l��c�/���|�O�����r*d���@�~��
dԍ�����h���̬���t�����3@�z�g�1�7�d�&�"o	Q�����v�=T����]U&�CMG)n��͆g���,����k@л,���M҇§ʍ ��+��o�L"�3������5 ���mn���!k�Ec�v�fV�4���/3�J7S7�~X�]h���?�Zj���Ju�n�:�R�6)��/'�mʲe��8��R�5�����O��U�%Z����~�RMW[�k�����n
ɝ���P�i��k��'Y��B������h�2���vhZ!�9�`lcq��9v�Z�V���~{����F͛k���8|�0��]��H*f��W���4t�+��	�;7I�{ER��ꛗ�R5���&-�����e�~ys�ڭ��P�U��M�e�I��V���}I�N�ѱ�KT�7j�Tc�%�w&:�ʨ!��8�#%:�����E<���_i�\8|-�@q7/v �$K�sI*3�?��2k�iP�T�m�BXO�njj|�-�?�z��.�7��Wa�i�so�u�n��@���`o��!9� Kl�=��ul/5吾���}��`v�^OK�ow$�ߕ�%�1qϛ���8��/_�7��7�^�L��x��΅{��zɖ�O�7�P\]s��u�V���;O4�z�%��fs��5[U#`��IĹ�Rzn�]R���a:����؝���9,M�j��i�Լ�P���t�e�˕���Eh���_κ_r���iZ?�4W�S���-3=�$dq�<3@���ΎӅ
�d�OG>��Z�&�:�z�+p�o��5�X���/Z%-z=q?��nq����DZ��B7�����G֙�6e+�@���j�z196��"P�B�����wm�a/�g3̮����g9�y��#.?3lrr^>��f���o �fWlDp��+����h�����L�%�n��:��%aNE	������j�(�D#������y$�1`"���7 ���>~�����)6�bnBo��/������bo!~��F�@7��z�wb�]�ٷ�ub����E��m�^lR'�,)�lr�� P�N7*b}�]�������[�	�E8 |�RL�,L���Q�,�bl��d�I����2å9�˲u4��� �-��C薕�p� ���r�1�}ʆ����ɢ���s�B��V�	���A$�$�q1����z1/ďQ��g ��h&H�ϐ�{����
��L�^D3����<��wǘw��e&��@v7aB�x��m��s���D���ٻ�O^�|[d�!�Z2|7BD;����V��|3\��#�F%'�u�8-k`]�e��ߕ�.>8��aN��1���xW�}7����*6�
U�P)�s*�1��58�+����ŨSŖ���QF"G٭<r	V��2#s��)ݰ�����[L��s�3��?����������m��!Q�h�$�r����<�������sT7���5��Ow�I|Ş�s�L%�w⣖���T��cf�x�3��+�<~_UZ)�_�/�zt�b���|�X���tѯ�i�h9���n����0������>��v���,�\�g���h�qT�mwo����=3��^�3��c��/Z�mS�mk��Ź��z����9=\c��+�q��
$4���Z� �ɭ�0�>�4� ,��)�Z-��@yv��|�n荎���4`�"�,�ħ��tɸ���Ġ�����M."��m����m��}��f2��o��>����P�g�鬪�.-z��t��~ΞO�Y�)��sH�x������d��T�<�x@�^Ui|�V��	ź�ȗFQ���3�t�@��ނYk���}[z(���k���M�zw�3�B��r�j�ܧ;�lw���sY�!N}ƭxʮV�R��:����e�Ta̻V��e��.i|�p#����s �f�dd��*&w�!Mg���l����}��T<��:d�%x?d�K�.��8/7��|��g}��g�\�6��Xq]K�5i��7T0�Ҟ+t�`Q�m�9����g3�� Y���n���A���{J>).���i�7ދ���C�;V�>X� v������Z�D[) q���w<�wy��52�]wf~����;��qVg�t��Z_�$����k�V[��1u�@�H�y���c+�����Ob��%B�wg�jΈ|UtY��t��D({=�	V���P�?k������u������1�X�[	���W3��
�O�<����4QRƵ�e�R@}�>�&��c7����X/
�H�*��C)F��Ύ�Lc��l�y>��"�n����t�a%\����x���ݮ�ݻ��5�Q�7�ݽ��<�}apf���>^��>����'/��s�|%��2O�߄[Xrd�a�7���K �I�;�`��y���x	���r�<M�p��2պЄGiP<�PP��T�Xj������Z�9�Vw��=J�y]��y-V�*����ur_�8)2���b7�D����\O��̹�w���PV�3�?#�bq�
X:��-����Q�ﻗŭ�ϚBݤ׃/.w�ݓ���e�1j�)X����vu�I�5%~�l�@���I��?��5t�j|@بa�8�@A�0��Jش�Vl ~�5���.���C�F��>�`-��Y�eߟn�cpf��>X&a��i��Ic�^�Y�]��T@=���	'�<����P;_x�L��lh8͋o����k�����Yj��e.�x���q��բ���& V��9�<hI�����M6�������i0�o���E�[8����=O��cz��C����v��j�"]O�<5
�\��(��B���dOJ�
4�0r�~�0i�����xi�C%^�U9>��/�^�Y��kٺ��H�%�A�)zuw[�C=�7`�=��;�eP=ja/�G�Ul��T"�iR��c
��TV���r�g%��s!��p�%�t0��d$��°�����-�d�*�������=��uu�H�&��P?w�t��6�kT�?@��R�vDH�{������8���9��冷�:m\(�@�?4�--�љ:Gg��ۍY�Q ���|��e�%ȮY�$%7K5�Q��Ke����ʙ���v< ;�ɸ�'�{s�!�P`����Ϋ��C�^�Ul�ԔO����2���*R�:���"����o@J�����Gg�n�U�Z4�%�v�жLͽ�O�SN�~ҡ��b��\r��ʈt��n�����d�UX���&�NX���w��T��b2T�X�Q?R�"�J9{AL^}�@�nfo���'/�σ�MM���/D�]G�qV�{��������\9�3��g ���U��gs(��Q��	X؈�k^tM����K�a:[`}\�c"p�^.�b��(%&ġЪu
��nO�7a��u�Z:�[mR�$�F���軄蝚��f�� ���:g;��	���P�]�J��z��橽-��_nSX��0��%P�,
'��پ�K��#�ًE��Bx"�"`X�(���?
����wy͞��%�[��fQ��I����n�nX�G�#�&/�?�n�=����#t[˔���U�M�AY�c@�+��U(B��P�d�t�g7��LC�����TvY�!��B�SҘ�F@��}���5�o��\�͘y�P�D�� Ƿ�`��+�[7|~$�NXظ;�߲� �*�G�>z ����("��.�k؉p��-����*���t����ށC�v<ē6TC��s'�IND xѠ����h�q �WI9�y�ݦ�E_P��l�U�i�Z���&;�(�"X@F3F�I�s�2����ݕC}{�.yu��"�ɍz}}�<q���s�֫L7��n�P�����s�W�5�R������^�ON6���B��1'�U2ӻ���-,�����^�7d�$�R9�w��{|�9!Sro��/z�H�Vi��E�*�ȣTf�d�<���� <@`�I��?ΰs�>�f'�
������v"E��D,�)|mU�����T��S��]rG,����7�e�N�d�,���EK�;�����-ܑ)��q�/�_ƛ�a(fŷ���4��g��҇?&-�b��$!}�Y�����!�	E�@j! ��٣LۊB���FJ��$�:(5D��lm�ƍ�X���bĘ�N���b@8��>�d{��!�^-W��!9��i1���ы�C�)�^B��}�:}P�
��X�+�J��.ƹ_d�D�/��{`����֙����	�.ŴIh�ZD>j*�����7-��$:đ_l6،X� �S�R�N)��	��{m���}�Hbaьߣ�-��ߪYF/��Lah�(�>iH�R椂��x�����5I"��.;P����r�e~�%`�i�~��4	����R�k*+�&��~g�_w�@��%���p��c ���lZ��K���{�Dgl��q႕C� �T`��^�����@E��,7�\��o]g>�K�?fF�8��2g�]h�`��{,��P��:8h��ijzZ�	���=.�v�5�	�E(T�C���j�MqZ��j��̞7�4�X��P����ooX٬�;�IA���M7��g���O��'��4(]�14�h� 9,�ssT��;I6j͢M���IN��kL!��2HTJ�1g�l��ʋ��kb2�K��ސ�[w�])R�d-�J���-��uޮ�"w�;�c�:��[��:��%��ݭ���D������I�<�F�)NՆ��EJ���(�����X���|�]J����i��Dr	։;��ðc�YS�P%|��әX�Oi��������������F�1U�|fծA�H&}{�eF��9��� �i��(��s���4�ޯH����[_��/B��9S�Oʲ[��8�E+�$�IH�N�u��lnW����*#���pΖ��6�K�����#�ࣦĀ��v*ƽJ�e�<Hz�����"qmw^�� .9���ΦU�m ���a�n?�| ���o4ܾ߲��d2�Ñ��qc�eb�~ā�I���XQFl�qB� 
5������8�^n�~�Z��"�*2�%��a�*��ׯ�����zG9��rj�dA�I����j�ì���ү��?㴺�H�d��rl��!�@^�}�ZL��a9�B�n�������, Q[�S?�>�P�Pc �f�>���N#z�$݄H��L�|�	��?���,m�[;.u�b[���ٸTߠ��I�,(��]3AҾq��NW-PTh��e��ϱ&��ND͔Џo��ޖ"�B�b�WF\�1X����u>���/ƹ�k��R��M�,�c���[�p܌e�]���¬���y�U����sX����|��T���G��*U)&N�*���,fFG����X�|_h��� O���l���qGD�x�U��X�
�6�u���t-O.�c<L��)�@k�������S�k�j�Lv�CC��j�uN�BU<�$�/�����`]��DܷVLC��9[0�h�;2���g��l��5�@�NO/.^N�D=~��t6�dO��0Cߗ��R0�����/��! w��i@��d�
z��b�j�z.?�A;��%�l���ޯ��aV�}Чښ }�Grُߍ}}�,8�=m��=��K����no]�\[�>"�lw?]d�о�ߨ�:E�\8�$s�p����<ii:K��^ �������3'����o�p���D�}�)?�|9��'^�d�1X�[x��Oo��R{��@#����7)��8�D�t����i�d�	����2v[�ݩ��=����R7��Q޿�Wxn����򽟢�QӍ�P���V�S2�P��H�G��J=	]��i5{��!l
�x�$pu�7�䊘iE��n��M_-!3xGL�{��6{x�~�����s����MmeP�ɤ�n�6����k!�X��JfEd&����k�2� ��
����٥��C).۔�����?��خ�#T����I�E�&w7�H�
�i��:�����o,X��`�\H�9�'S��$��
p-04���j$
��ݚ�f{P�E���W�{:�w���F ��#Ce�M��0�^�8�~�p�F��)_E�S�H��t���ws���R쎭�������X:���vPyoM~���XR�Mҡ�޺���uFF�V��D�ѯk��Ѳy�~J����.]��.�S�s8�hɃ��ǲu]g�"*kw&�s���!�E��| Lt�Z��<� ��Ώ�FEm����c���_�M���|������z�#(Æ��'��jݐ޲�]K�e��i��<�C��h�h���X �+D�V`i?���:~ �O��*���7��V�v8-�煮2$���ݟ��L�� h�x�$J,.��4�"7�mȻ��D�?5�Q���HSr��T B�ݣ6�X��	:΂�5}���`!s��v gʤm�m�����L!�\������7J��o�X\�b��2�L�bi�%R�Z��f�^�/�D��jTL��>��S5d;���|��G��ES޸�D���J�۷�)�P���%�bI�p>�`մک�
#��I�8	�	�ЄQ��OJ�Y�,�/�4�
��f%�k��y�Z/��A�O�'~}��8��ڸ��
B�G��}T���~Ҹ(��FJ���5xx;g,@� ?����T�=�q��n�1z&"�#Ч1P��W>M�/�P�Ӱ�)�3-H�G�uf��)<�c{
Ghf:��ȿi��ٶ���K�:O��Y��'�)Dq�0N�=�E�?	�%��D�؟�����h5�xBj��	�*[T������XS���{�(���j ���}���sp�WM��� ��<�����t+��)`�I����1��|̧##�ܬ�����|�$2oI�L���L=Bg*@̮�q�O�Ty��*_(9=g/d_?�E;�/��LZ�����z��LH�]p�^v#>�2o�`�x�Fo��hD�ڴ�?F�m�v�%���"���7�s�
DJ��W�f��~�FR���$o�J$�7B�D�Q����*@�%�g	f8��w�`�1h���TNf�.��[� ~��ӡ�� �J��<��0R0�bS�z
7���n��e&$t�T�Oӄ��P���3-*pb��En�ju�t$$0f�M�I�mS��3�3���-D����2�t�p ��t���9�v�@U��9̯ˮ�%Bd� �M�!a�4��P'�ר���s���9> }	*���E3"LO��(g8]܅���������2l����!�5^�Ϝ��R{y��s����Nɖ^�M�t@q���Ĺ�d#�T��ƻ�c���0�obBჯ�~{�����.;Ӡ�;2O,l�ʐ����������"�xc]')�U�cu�,��bت�v���gia��>&ٳ@�����a�AB��}.�'��p}.fg>�3L���O�u���/ �&��;ޞ��V���q��U�f��-my���$t���b�3��t7�j��#����M����&!����1Н�TV��1����K�`7�=��T>L���9t��'e
���B��A���2���Pv>����I�,`�� #2�D����#�z���&�^�-]��|����O����gu��ch%�.��1�\]�$�\�e�ZN���υ�q���ۻ�d�*�n<m�1Q"Q�#��u5_K����:3!��Uy}eO	�ӯ5 xՁ�M����=]1�9j�@n%$�M]��ɽG����7�&1a�Qg&�x�%�.F�NRu4�yqI�\3�c�-� ��t��6�`ǫ�
0�ÿ���n6a�b�@}$W�W�f�AY�$��N 	��CJ"��/5���
���!MSѻ�W!�� @�F��:��|�[���|2զ�6f���]r���i�D�'w��fe�K�����^��-�!�βȁ B�\��*r�ut�fZ� �b���ں4*���(j<��N��P�&g r�JT[���g�����B>����tk�L����>Zo����0Cݓ�. ��-��`a(4�����T�C�Sg#_�6�e2i%��t�Q
��haS�Z�G1�5_Gr9�k��+==�O��]'l6�@�o�ıN��i�ݍ��1�m���8b�P ǩ�����
ÿ�O���`�����`H�Q��&���~�*�;���O�8H:ȁ�7_�~�+���8̆:�!'���Y�q��t�dT^���+<yk��Q`���=�v~��Ab�U��}���A�6���RlbH�{��=���ٱB�J&����ן'�v�9A÷��,�� ��~�z'p7gw���h��\)�7k��+��'���%��J�	�|�L���6�9�� O���~ޝ(JG�El	Xr���QYP�a�R.��#ϸq��D�h�mk���7��R�]�Ӓ[*�7ϑD��R[@���1�F`����9Ӎb1q�"�F$8<��
]
���EU!o����8�w���UN��i���8����Ɩ駞�M����+����:yP�4�����UX��1gŋ��_ix\haU���X9� ��z@3�޼H?���c �M��GAz,FM�KDBP�9T�w��8!J�jf(e��
:��u�XRrS�I'@��۔�6$鐇5�a�k`7����o�tmJ*Qd�u�b�EdKB`K=���` ��wY�����Tp[��;(b*����{'k��	��L�B����"|^G��.��
�C���Z����&��;PVVI�%��?ݶ���yaf�"DU�Q/�84aX�Ab��E�����yE�@��Fd��A�	����"�bl;K���b|�'�6�	h\��E�@��Xd~�\b�Yk�����z�,6��~Ŏ�柃 ��m"
�
�;���y���`� ��ʆi����K�D�"f�k��}��Od���a�9Q9��P�X������{$�O.�,����k�j
M#���(@�_�R���>����a܃V�������O2��	�͡����] �� ��Z�rXʿm�.a��DiN�e�v��anԑ��M\&��|`Q{_�*p�`���'Y�+��-�H�f�Ɠ�uC�II�� (G=�<�0%�/�j��f��e�������P^cc��_�V�{�.:�G�n~��Zq�8��?����re��%`�5D��`A�s�f��O�cAfE� e���f�9P�᣽3�5߀Vq�ƾ��4�EϺ��������D�]��;M`F�n@>0ǂf�4|�o]��*�2�L$��ɽ�rr4�>&{Q��_�qp6�y�`��D�F�~�NGJ:�E%$m�.��F���2_>�+	͟L�o��qU�J���D�h�2;z"��� �7�L��z|�G+�6�������x��D)%��b�I���Y
��o�'�������ƒ{��或/3� r	1U�h 2���=�7��=�Gu"��(so��J&���\|8a��������=�J�
2�w�)�j�`��\�Q[R@�`S|B4�����
�k��]��%��2��K4E� ��}�6K�F�J:M����>���k�6b<H�̩d��3Rg�����I���$]4�?'m���Ue	�Z}-����Q2?��cD��R������a����:I�-�֕����^��P�~`�V6"-N��ȸ�e�&�T6�t�
��%��vւ�i�`���xݾK��/K/���X���1������w"
���G��0�|�p��p��7g)�T{�\i�G�Ư�bc����8��Ѷ>bS�qc��!����_�=���s.٣©�*:�zK�"�ܽ�׋�o��elOq�������ҡ�򪝎\F�X"[�Tg�?B���pa6�2�b���Ŭrmn�O�
��Z��qHオ���',`�{?�0��]H[�:}dҿ�[��������9wu����wJy�8��=H�5�z��-h���=�3h�A���;ҽ�]DN��?	P���6l�[��a�;�xKɒGG�
��>9>th�yot!�T�`P`^��#{2����.P��n}8G���̌+�����MzW��9�4?�;K{�-�g$��+�y[!�Has���E||�_D�B�<o�I��C3.{���4b'��,�8��8Y]�|ʑ���~~���j��Ü�x�����0��Wh�xө��`IdXslL��v��t��Xn�j���Aȷ��=Db	o�ֽy�G��՘+��	a��DD^��1��W����~�3E��4���--[��X��bQ��u�����&��U�H{a23�
�P9��4S��i^�v�R�/dO�|#\�$�V{U����i�i4H��Q��hGS��@���<T}7%2=�eq� F�N�W�6�p�0u���+���og���pu�B,g���O������ XK��L�d�]�i�8�b�F��+Mu�W�6`��h�֯�Y�!_��\>�͝���I��o��Al�_PI��xK���3퇂;
�� ���z�Ņ����G:2�H��d.z�D�4 ��W�
2�̭�S���z�e��Ce�����1h��q��ۍ��u9�N����N�������+��o��`#�m��3P֍eNI�`*��䊾09C�U��ŷ ��u�2[�f�l�3���[x�ԃp=���{�.�e׵-�|���Y�!��e����]�'���=:�`:���5����k��V:�5{���*F���t-`��eaY�*n"��"jkw*�Cֿ��^�d�<A�Hw�&)*}�_.^�j��PD���c� �hj��?�F�܄ݱ��S4wʤ�k�m���<��r,���>J�ƀ�����:5��؂��:��}%��Q��r�ޱ-�cNB����6��_����b�O����&,%�fl?�v|e=c'(j�^k5%���DϬ�ܣC�r�M���!#L���z�3��a��a��!`�m�L�R��v�l[hZ�ÌB	y���vwC��(�����=�.i{���v\!W����u9��jPX�cw�OY�w'��}��V���#� ��;۵3��J���ɤ�T�M6�mA�F�ֵߗ�v@�I-�f��b�2����z���M!Z������y��Z�1X�`K(�Z�0�@�w��-V��d)�<H�ӧ�(ں�v����'{Oמ�Z�n��1��V�a3�#�l�;{��kO>oѳ-���;}enh`���Ə�1��k���K�t@Q ��sx�~���C(�`k��
ZS�k� �$d8��S\4�J
{���=q���Au�L�X�]�$��þ_���44Jy�a^��b�IQ�-\��&����RnP�eNh0�~��RH6I�x+U��b�\*�@��K�9��!I5�o����R(v�J:)��\�v_g��Kh,$��R��+O"[����#�`j[E,
}3;IE� 7�*�6S�i��]���
��W;�N��R[U�lQU�_���8T��pngq�:]KD���"�?z�6.kW��T��&q�אۻ��.=�4n�C~�)
��DB?VU�n�m$G"��u�2=�LQV�gh�N �g�B<�����ˇ��9�z̭;!*���SvIp�V��Is}��g�.�nJ����U�F�`�<㞢sU�����)�S�(u'�c�H��A�K�h�B8*	j�z�	z�
'���u��
�ỵ�V�:�DI������p�'���s8�b@��	v�u�ťKҚ����V������=C�-e��N�-���}<F���-�>4tp��-`�[n8�c��_M�	v2;y�D�,-b���)2Uz�rn_K@8
t_R\�_��8���+�`��`&1]����g,D���o�<��%Q�9�%7�%Go��$3zk�c��奊Y�R�� ���I]N�H�M@��זn�_K��{Ҭ�/����[0��;�G�-m�~%�P���J;Sݟo�wP)u8ϥ�z��l��0ɜT�`}?�FUG�8�=�\Г��C�~3���>纁�a#�Dyu�e7���d���j��\=Tf�&��K�SZ�Ɏ`���a�"��P��'45A%Yۘp��Bo��N�f
��ն�^%[����wk@���Y����q��ѥ'e;��^��6]jq�g{ 8���‐S�&��%�5	��fʌ�X�d�������UK��CI4�îvẀ�	%lKݯP��D-P��Wf����GZ�˖%�=g��%�-��Xr{�^hK�VI͇����G-I+�_��8�Pj�0t�~ �m^�D䱯.�?�XN�U	��'��i4g��Q���c��j���ޔH=��]��^5D\�A�K@s
��-�n@^��
�2�[�:9snu!8�T���(�����H?H�v37P�a�{�3���z�*StT� "훽8'H���:�mqE�^j*{l��&�'���a4�A���7^^I�����`멜S>����f{��{�٘v�ZZ�Ǎq��L^ۮ��g?��I9�i9 ������o�om��`G��\�������b3�)q��u«NBP�:�d�6 Zo�*%���wڤ�&��&���ý�8�j�+wl����N$<�%����-/J��"��}��'�g��Y��~����!�$3�k����u�5&�t`�&��V �z���\����~
X�B��Pv@p���N��lS����.�k�\X2��U̫h��5�~�|?��o��7�b�^)c?oX�W��}�G<�U, ��l� �;�����$���Í�0��*7���;�L�9��N���t8��w��^M�����Y���]�f���z�AS��֑���W�b}��� (��@�:��La<c ���vo�a���i��L|�Ui�1c�`r9�1�5el[�I�s�a�U"���#w
�qP��
��6�2��du?h�S�A�
w���� ,����MtH`�; t�K���D<���3���׊��N0�-O��$��\fwH��P�B�'�Ã�f
���P+Y����s������-Q�K���@y���(�!H��L��uA�|�NuŦ���p_�rX	��U��n	�� ��WP&����m�@�a�������@�;W_,�zt�7��7������a���O����;�% r�O���Ђ��\���,�G��4^c/
�R�-S�� \J��vY�i�$P�Z�w�N��S|�BTD>mP���pT���\</���M
��qD%ᮬg�C�s�Ⲫ5=�n��u��E��M�M��g�M���v��b��x�2s�M�}�
��vGi�KRa}����;���M�G�Ѿ�<��Wjȸu�� t?h$�;πK��)�g�_!���=^Y���ֳ;B.�Ly����7�����f� ⍭)�����D�w݁���k�� �ۺ/Ht|^oC�t���򕌻{��{�VZ�~�e�)06w��z������fD�)�ϑ&�B*���x�#����������uW�4�mP����h�ڈʔՍ�������O��1?�@��m�����Oqۣg7:T)��������K
��ʮp�ܚ1O���M,���˹��Dn.���!]W�Ө�G%���:,��Jl]d"��Q����<���j��B�<��`x�PZV��f�� �IW�����ӂƵ������zt뿤�%}�uS{���Z?�݈NRQ�H�����b��&�W��Tb���|�dܭ�;�;�qU,�VPK�^������S'@�֎J�%�l����/�m bbQw�넧�ϭ�~ᇽ�-���X�_T�Ӵ�i$��RǛXLд����,Qx2z��-^��?����_���Uۍ�h$��.�I:js-?:>Ls�J�y�h��+x��6q��b�?�K��$�
ťTk��\R��:P��č�pX~��V����f�D��F=<H2�ۅH�L5=���n9f�eS��B76s��i�-��X��[B�����bs���u�x�c��nm�,����V�]����영Nb��1�ZŃ}9��ڟG 󵚥���0ԩぴy&����?k&1��?U�}����Z_��v�������L��'�嬔dHf3>nv�^%�Md�2�2}��4��p9�x/��q�eg1Ym�YX�=2����qb܏%��*�KCCu�&�9쏉�� �ۤrG�H�+���-�(}w㒪��Ĳ���Q	v`ij[^�g]�� d�y�o&�����ub�W)�%J���2s����)z��s�*�S0��W�<3�����\`Kw��q�J\F����]�o�ג���Yų��뻇��w]l�~7ch���$\cB��W@A	��K��f�3��r���yKMR��=�Zu�E��v�C��{��幞���>;�X-*��Hz*��r'�o���287��g顿�����p[��IM�+�!�;#i�%��,E��I�����j���s�6�w�;�{,��}�������?�e-�y�n�dp���#�Թ��jb�OW����w`-Q�j[	�S�e)��Ph��s�A�s�W���z������u����\a�ҙ��K+�J$y��M�~E���'�`����3��Y5�լ+�w��;1�� $�ق�p�]���ݽ��fC\#���Ϲ
(���+Tևڥ�w���'/a���iR����]���V<P���{?�7+��aVs�׼�$}����Yw�m=a<�L|���>���*(�g��<d���^k܄��{-llE�U>�GLR�� z%9;P'z�G�YF�S�n[#�d����]��׍V��`Q&�[}[����s����9i�Ѷ=f핽����4�q��������33�xC��Ps���o�ՎZi�حng�q�d+�&ƀ����LU��]����d�T��!�)��fef~R3X���-TGo��8�=ʇT�G��tn��O-x�B�r|�m'���DHٔifpG�rf�Í�π5�qv{I�!J�9T��KE�\��+�k+Ʃ��O%+b�
���q[�r�xB�\z�_π��1�T>+U�D�� ���J���i���Nm�jo��m?Iqg�, O\���ki��!�~j#�>0A}��u.�|��ĝsS��T���	�;Ol���I�/0燛��E������x��7�so��[��VTJJ��P2��m�PIȘB�1dO?E7�.�2V�̉�1���J(2�$�1�޵�^�{?���������g}���}�����*_�� 3���v'�˘�Ï@��}}1�����[o	w�ybG>
�+��z���2FTCދ0c�����6>{� s;|�{d���*+]�ٝH�]��<i0E���~��F��Č����fOl;�����%�ڿ13,�㬿�(.MƖ ���>KH���0ad�J%����B�녧�~ �o}k�7�_;-r��O�nJ��b�v��`����|�P`:a,� �x��Ir4��,Y����%Z�N}}��B��r�O7 X�Z����IL,#X4���6|��U��f��	�7��iH2$�lqX��K�"��%�STJ���T�+�뛋ϸ���V;b-���%�j�~t(,�B�������v	Pw)�BUװ��i�S�!�Yl�;����e���R4�G�s����R&���A��)�"S\�	�;��T����mT@Hqi�y�ga��:��&��,�z�
�zJ^���{tF�
<�?��"��/gO����w��xU�Y��#�bi����^�84�+����~Ք}(�O���@���ҹ�͏bJ�re�UJ/�q��8��w�H5 c%�8��	�u44��Xu��!#\QRH�8٣�̕Zc��S%��|�ٗg	��p�p=��1��롊J2�}�Gkp�N���O3�l�T�ʴ<'<Ɩ��6$��'x�pUZ�<���Aȹ�|�f�����E��s2k�H�R#@R��A��S���ւ��[��\��Kq$���)�����xH�uvV֠U)b����k�7r��[ ��S�>1렔}�ίn�8���= ��U0$�w����"���*7� t��v���O* .��7��N�8g,��7R��̯?�A���c	t �"u^\U�ʲ׽��w&�rIي��^O�[��m��.�j0�V�m���圣���,�7�4~8��~RS��'A�tv)�J�; �Ȉ}�>Tx���{�z���p�n�b2������V)��V)8L�m[eoo�G��KJD�?�v��5?��˫�I?��R|�#�����Τ�?i����+#�{)�t��/L%<8C��Ɲ�/��6k#5�4v�2q
=���l�uo�/L9�b[e�����̯z�ƀG��Є����d�NԸ[��6�Wӧ���{[�L���5�n�1�U6 V�|p�X�⾆���Θ�#������D�#�p�O<����5�E|1~��ͱ+�7�^?�EX/��ǿ�U�-�4-��0�aS3�@��ӧ�+�$�
e�I����U'�U!jqj]2nݭ�m#+�����c�4�Fs���ރ���e�$��^�x9��*UF�韍����Mw35�,U��r$����)-�Y�p#���{�u�K�,t5>�M[����^ԑ�{��a�z��N5���s���x5�q�><��68/��E��F?�oߦ�	�Ur]�}�\�UO_E5X�-Y�f����}Ʌ~���J bo��(��DD�7�뢈m
#3'y�B�J�I�9C��Dr�l�s^�0棹�{U��0�wDzM��� �< ������u����v;旳oߴ��vϖGj��=v_�����NKň���$oϗÐ �ג.���!R7D� C��ex�ǿa�p��z��yfr�*���`k�}V��N������Gtoh���-`���%�N/���4��_��K��/�^.s�耕���%��hu�I�X��nL�u���g�6�R,�>�{԰�.�1�;�4�d�Q�]:�0?��� #u�_�v��m�I/~��DaER]%�A.��υj�O�ֲK�>s�ݛUU������77�Ϥ�uț�?'��<
�j� ���%�G��]���t.��ːܮ�^�fߛu����ԩ]�!��~QI/Ĵ"�ވ;Ʒ�rD��\|G�V����?_V~�w5(���k	���_����c�����������~�ߏ���?�����~�z���F��ܲ��}5����{�	x�?��d<F���"Աd������QgϜ�����=Q7r_'����^k��b@��]Zk3$�m���`PǨ��$��B�4_Y;$��,MS��rjω+{&�"�M$��c/i�y��D�vy���oX��b)>�48b��k꽋Pӂϻz'+8��/���z̎��>\���Q���?�Y,H��@VBM�A�⧭wE��L���O��61�;��sF*<2�\���.��,��#�5N9S{F0#L��O�ч����|�9!���_[(C�;f~o���X��͏.���`���7�@�{~#��M��kpKt�u����Tǵ��Ϩ�*�^��DiE�%y��fGJ�-�6~�&r����=ﱥț��r�����,�y���;�	2��������71	�\hLa�/��&.�>Pݑh_*r��m�M)��k^���"rY�J������-bm\�������hB����\TQ.fJ���ٴ�/]�2�/�_�W��v�\���C{|+��R�H��ZΔ�������zXLaޱj�?<�s���/)��X�}ؓ����	^̮rQf��k	�����}�/<�4�i����_���B7�j�0)�Oo���/A�af4^|����욯ƕ��W�8���Q��U�r�]�{�U���Tj�8W�>�^�]�Z��p�3��?�͸�9vL��#h�-u2�W�
m��l��G�fv�;�\lx�O�o�L�������W��G����n$�F5��qa���W6�J�:��m�ae��t���u�r�� 0�8�t��s�^L��@l��u�u�:��.�&7�z��A��a��/�z����h��܌n�>�!���eei"5��C��[3dQ�`��o/���2�X���g�]�2\���N�;`�5��Sȓ+PL�cT�G{G���2+i��d�`�������?.�W}�f��(�b��r���Ć����.�	�����5r�~�ƭ��T��]#��:u1��Z������+wjB�L��].v)%=�&�C;8�U�e>tG/|e�Qs�rًS�T=\>��Z<�"����/�4j�"���Z��t���S<�%#�D��q�j��>]���Z�A��'�C��%�h���(�����$kQ��� �D���&�~�`��&-]#��\HG���l�[��4��Ы7a�o��m+!�x�Ջ��N�&����4h��Q�"��j�W9_�ӶR;a.�Y��ġnZok��W]nl 
#_��%�fT@SUw{���e���*x�gZ(�f����
f�e��5-��?�I��L䉔5z�����fx�R�KZ����x�)l��5���� 
�WjS{a�_�O���ܛ�;���S{�#�qD͞į�I5oe��r3�֪���8�l�]�cba+���B?XM�'f�vLˉD�0̅[�9�]58/K�ay�E���,�j�U���f@��Q�-?Ř+ze�6��q[�?|��/R5���EC�/��-��� �2� C|JBw=����vls6��$��԰<x�.E`��I	�}`4ou9#�ί��o\�K̼��D��'�m�X���&#��8��C^N~f{�\��Q�,	m�}-ݮ��=��z�T޲��$["�=�r���Z+���y��%��Cͽ�-Z�J��Iz��ݦ�H��%�ư��.�8����e�l9��"sS nQ�i�Bw�h�ё����㱘�_?���P���q�� �o��iZU��rގ��n±`� �o��Py_R�9�'|<��@D�	����O�����r�'�6Pِ��ˌ��n6�ij*7�7lpBȾC�ø?L�:O~�8�r&	Rzb�q};hԝ��bq6E��K����7�f���n���E�4Ʃ�FQVsaL�t�v|�j8=� t�q-3����m�h���N�\�z�\���t���7Y�����6�Ӵ
��@1�NO^�|ޝX����a�Y	�/���] �M���	��w���7��5��6�¿�9��o��7���ݒ�1��uMQ7^��^������/�in�>��>�Z�?�^���0�}P�n������/�����)R����m��k�6����H��<\�� ���x}{E�iL �XP�9ܥ�S�:��w�V>c��BU��7-_��Y�ϧ�ǅ���? y����~�� E�;�6@/Tyf=�?:Tje\��������謊�$��<�Ǭ��������G�Sc??Q�6���?B`�C�D��pg���q2l��.�~��2���%��{h�(4JB��(�{YF����J/S����r��w�@]��z��1]]�\��1g��h�e��Bb��փ�!��?/�v^�6��i�A�[�V����/5�0+o���v������gJ��W�B���N�8+���(S"�s|_0��+W��g����n�z9g⫓�Q�~ʄs��d{MB�-\��B��K�MW<�U�b�Ɓ/a��{�D�h�iQr����b��\�B�\�B$���D1��Q�� N��et_.1���_Hjۮ�3�zq:�]��l�v���xܷ͋(B�r�����,d|�A�T����emw�B#��8��!SGm�U%��R�#�8��)����q[�S�n�-�.��\��[s��ͭb�& �ҍa�5쩢B��1�}�\dzx����������&�·���ޑ���Z���1|͋1��2U�!f��)�����G{"�����DP��;��!�~V�eum|'��4�3�%\���co?;�Z���Y!�;�t p;p������O�!�

3}�P�n����/WU�E�i.(��n� �J�c$��Z��Z,�mw?�A�j�<���r�\�ǂ�NݵP���bx�j��v2�N�*�����0��:����d���@���j��.������󮓍7���Є�>�I{�r�g��q�&��K�}�m㋑0��6�Y]�^^sã�% ���<ئf����!�#P̓]!�%5�d	��B0�bDA�g�E5�=[�۶m����G0A��HO�P��'�O���e@��<��&j\/��#L6Z�h�vt:�#+�o*Y��ǣ�>��ͷ�5]�A����]�75�r5]�#<7>Xδ���	���mkZz�o��&��w�XZV��K�D������8���P��D��ti��RU�d�gM������z��W�d&�)]�N�_�O�"�ޞn�T�*������A���8���]Z3SF+�~�-�p��6S��S��^@�1�w�?�]Z�YPu��3?oR{���'�i�ԏ��m-�:�:���Q�����,����e�J'R]�^���s�"���PI�x`�o�S��	�\�I��eX��)�(y�}��#�Ȧ�Ar���.��$O4�w��"b7\#�����u��G�bXWi3���IQo:�r�c�b��1�84=�H�r�[�#p��e�� ��3�{ŃF�1�]f��� ��KD����Q^+;��9�~��&�U.�W�b�\��0�M�%�z��X�;u���p�惤��MZn�Q�2�ۤ�t���4��!>�pi���vm�MѰ��@�m�okT������y�>&��%�1A[ZA����v��qW�����6ǽ�d�H8s�NT���J6W�+w��1�R�d{:�$9���x�K��/8��ZV��{��Ymz&]'�sk�Lȁ��������t�t`Ya9��1c�<�a�*� ��M�-���sig��Ʒ�Ąw9;��H7�]�=YI���t�E?���J+��׼�r�ϟ,�t1�J�	ty�_ENI��z�x0�Ct>մE�,�P��i�["��xX?I���d�`��6_�������K�������?��1�b;Y_��6�okoh����oQ^�V`����1��e���Ԫ[��]%vXhCy��z�{@�l�ʹNUb���K�p�����oZ�E�Z�f�V�n���+�J)������
6�sl�8�㻣�l&�쉣�!gC���q:��W?��0V5�W������E"7+����
�Cb� ���,�9mR�[���ݲ{�o�7e�^�ͤ�(��d��!_/N�&׬c�&٦��3�*�M&Q�'l������C�w�n�TG��1q��5���DM�y��5f0i�� ׳��1�,���Q�
�_��4�F���~c����\����6>;m�i���6Fo�SC��	I������yե0�`���;��4=���HЀ��9�#1���/!�w=��`{.��n &*�/��U2���Ӱ3ig7b��گXb�bc�����V���%{�cD,8#>	|�(Ӏ��՘r��aʟk���4�n��s���C�Z��1�ˣt��S:zl|t�m���ʵ>�@ڐЦ���M�P�7������{�m�ct���>B�%�ٴ�.g��h� ޔ�ؼl[}����2�0e�O��fw�ϥ����9� cV�E&�>�x�-nߍׅ�h%�
 ��a�ܬ�E/���Maʒcv`yG�-'�`�Lq�̮1yU�<$���&o�(�΅�� ���-��$�%�N%G9'C�`-������Y��.��ECp������8����U�?��nw��d��
�����Jx�C�{B��e6>xTM�/��߾�0�M��p�K�Ʀ���n� o>�ax�~��ݔb����=����<�� ؼQO��=+qs�Yk%hg�R�����l,S�b��o�U�<\����o��S��ȟ��M�-hq�l��ܴLL�R��X�][A���B+<�����Vc��5�,��h۝`#i_T���AGK��Vt��}��{�rtDBR�$;%��衏��� �a�5ϛӼ��j�;��;�abp�A�V���~�������-��	L��Z]%^/Z�\�*��Z�x�~M���y�@��1np���$���0%�5�������]���?'���f�%�7��z�ѳX�o�q�F���I�o@f϶�;�q VU�@��]��nPu_�@\�'WE/&���}�5ƃ�+pL��'�B��2�����r������;���N�a�&6Uq�{�m?�o{uDɳ�|���tzL��苨82+o�v�Baoz�`�@�� u�0���b��W�z��D���U���'"9�w�[ԫ�.Nq���di������d�2[�Nnƽ#,�̲*C1ꃄ�o��;�����0�'�݄��ԝ\`Ru�E7�m�"e#].�{[$�O�eMg�MQ?�Sv;\�j�dP������2�*y]�	Rɍ�Ó�	I�X��"�s?�7����o��F�v]�����y��}���fc?5�<K`�{�
�d�HӁ��e]�&A 1��#=�o	��(���`�3����Y��1�Y
4ܰw�T9_�H��ݍ10\����%vPo.an���D�NƃӍ���I�E��5Ly�!a�
rVL�^�Hvx��J%S�����)RHy�܌�����)q�}�"*�M������j*Y�?^�%�]�v~^� �~��i�P�V9�\�ĜxM�{;[�2Q2�Q�\ @R�^�e�g�U��jƱf�&�M���6nH�-��\�7㹊�$����ʲ��ɦ�b�=.��E�<1j��u}Co�E�X�����@��Et�7
C�4$�����u_�Z�&Z���	ZS�M�^��tQ;�Ά^ÿ��v�X���ޞ񂖋�$�Z3�ܰvv8r����'Ԏ���poJ��H��'.̺Be�����W�~5���>�H��\�d<H������� 8v#�AkH,o���D���#^����o`�O��Z�d�as��ôF5�ީ��.U� �vk`eBF]e�/?���7L9ɯEOQ2��]w�l�zE�%�MQW v�3��4�i�R���d
�e����[�p�|P��0���G��7�}���F;p�ob�ڍ�>%�V���ז��i;�ڇ�ə�%#ҬvH�����(>�v�l�O�f�{Q3��S�X++�� ���([2�����ؔ�Y��)���Z	U��٦�o���\^�p��p`��&���֍�2��:3%�V����Ԥ����!!���ۈ7C�e���F�����X��e8��f1d~핥s�J�i Jd6���(��L�C~�
�N�ץE�4���H���ca�$��8~�qri?�����<̚��1��K9ylh�)�&���h����O�*d�4��Yax�MC�
�mf �q��ݩ�;r��1�Hu���#�"��Q����KY�\�}%�}��.!xt+t�~6���!��-����J���.�Ƴ3�NTA\#�f�7:�����u�J6���8��纜��!����s�&��x?afDd�TFCN�#\ْ|�{���H���|����'jMO�5�Z+1�ؿe�j�Y}e�0nW�U��Ƌ�,�$�|�>�%�>�i#�>y)jn	�&��niN��iDhRX���� G.�����@tġ�G=./EqF��g,��*��ɍ@F/1�?W)/E4y��_C�0��w[��8���9��6�|-~��Z�EOh�*䔏�.�$:3$����C�$l�0[I�E�0�iI��n��Ʈxd'	�"3�k�h��ů�v����CMV���q-3g���	wbz�A|�8aj��KbX��2�=M\!�F�.p��pjA2b�(��FH�� M�~��k��^����%JJ� eС��[�)��5(S�mS�WZJJ�8���(���N4#ޜܾ���K�<��%`����Z+��#������`��3�af�zF�N��֋��q�,�[��H�Į�����bI7䮟FH�	C;���B%�4g����61D�Ǫ�w���clG$1ʼ}����&��\��d<r�A���!,�$$�F��ɷ7�v8X��:�E��ߚ1��U�*�!����]׀&�)�y<ćP2-�i�x('�GQu�F��w&&�0ٲ �t�e�����X,mKI��M�:��������'a���J]��(�8�O�-�+�o�����Z�R�/�`>d^#6;��+�]�|O|n�`��-��Er$��J��.:+������|b񚘿J��H�f�\H���b�r�J��]g���s�7+\ΦJZ�2e�oVR����7����`���c����c��ذP���Bt�n������~��n�C��G�v�N̦2mBp-} �����Ǳ/j � ��nݍ>�J�Ϙ��Q�j�!u_v}������ ���'�סX�)ȵ�M��O�N(>��j��e&�� ��e#+�ݴa�z���g�ŗ�Ѱ7Zg��2]@Ӥ��~���vπ!Dh$�'��3#�J]g���KV�H��ã��;�V^@MW`��3�5��~�	���x+����Ճ���X���(,��!�_����b�r}��Y�mr����d��-�F:�mA�Z�p���$yo���-QӢ~�`a�+?xǟ0 ���9�5P��j���y�a?�H=n x?|3_���rb%���e���`��\�#������G�f�24�$�a�ċᾀ,��pl�Q�j���"�v3�X�	����347��W�}�ي��s[��Ԛ��;�Q�XP�T�����cs{̴y	��:jqѳ5=^�rǁ��u��/w���p�����Ȍ� Pn!Z�7���W�يE�C�bEE�Ǽ�L#G�x��.=5�0�������%�~6먇����F�a9+ݼ>\ݓ���a��@eS�����<�2�Z�����¦cĳ �����q:'0h`���$�^�/ʼ���)��P��+��\��f>��-�*����̜s�H<�����'��`��"��^�S�1N�,"W7�E���`�	��X�2�*L�a�}���F�{�}��ZVe�_u=�
�g,���0�&��=e;��◗�P�H��3|�w��\�%
�bv�`J��^���`�2�A��֚�|�P�Ա:�a�8,
�]R:���&bUab�`]�ƶO�j-�=K1F���GB�qU#<�++E�*`pV��Q�5x�#dĵkq��p[	+�/ʮC%[T�˽QB���R���@�J	�ׇA��;�E	&��j�����6��H*8��Uݳ��<S��e��7��VĶJ-Ω��Aj�@�����5Q�tB�$c^t�@�hA��n�6���+���M��fk��(�H^�5��}C�l��7�� #�8���0rd.'ZF�K"��c$�����Lb��eՄ�E�� [a�k�}�}���z�x�|¤����1{�~���g?`�8���;�u"�> �q�N�0��t^��K���	B(��V�M�pR���I;:�j$9DO� ������xT�%Io��_䰼Z�xz��������)�E� ����\B�|	��" �@ ����7o�(I��g'y��6��m�1�vPe�\)�V��M�*H�Ы��z��^{oY 4�k���>��3��eYab�c9�����N拘���b��q��J:p	���wk�ܨ1D5�kw@��(��91%�z-/��F�Xo��1�>��5���F9�Zk`o�S��+<R�"ho�	?�
7,��Y�ȁ~'u��*r��
h�T����A��������h�+�^|S�D�e�W(�t�Q�0#�`q2�c��dNx�ؾ�x:�U�H��!Xh[ޛ��)r��~�I�`��2ў��
�jE7;�~��2��$o�ްP���f�|�S��w��
� �S���*̓>~���K,��2�&F�k@L�"������6Xc����ɲ`jڙ�G�'��D����ب41"X�6=��G%	ψ��`&��̤���/�"��&��v9�`����}B/� ��yQf"��6�7�����k�yyNs�]��G�n �\Zz�xO�'�yjl���
�'jί��Ѝ�cqF�Bl�;W:�ܛ@����b���F'��A�N�CkBq��8�Qö��0�ʒ�ѭ`ʅv���5|�>=�S$g8�a�&��=��>��S��퇸�1]|��M�X���ؠI��!XV7}���;D-i.qQF����wE��k�M1�oBya��}�
�c�BN�����̏�7��S��ߏ�W���}��V�|�W� CRl�j�V��'7�x�`uI�z��4*�Q����M�Y3�*,��B��Q��`��Լ��4Zz�ۤ�ˉOD��~Gt��eK��4�t�B(����]�o�rl�D�ƫ\M d��4��hg���!�_�@� ��i����G�e�ns��Ԉ�!�r��M*��t%1����;��J�O��J�:����M�w�/u̡�
f�Řo��_Ҟ4a��ꨍ���-��g��%h敿�̬�=��E&9 �� �JX����L��m�s�Kx��=�(��F� ��B2&���9W�ί�Κ�#ƃ7�m�>'3m6P�U�15?��`$_�mP����
��g�-[�"Ttb�t���+�����"C�k�1"��Y~_�'q�丶�7����F�<uv"5F�{HMx\�/u?_�l{�8��dXUk$��KG4w�q���j_@�/n������G���炣��w>�7�1����ݐ��V�jK�ܒ��Dy��sa��^em=eI��R����!�=+����+XV��췚[��q��l[h�4�䫊,�M*�o�[e�����{�ݟ'��Ow�GPuE�-%�)�,̝��EN�̰A;?���xJ�F�\qt����ϚL �J����o��a�NG�-a��c;�6�ǻ1������-�,�뺁1�F��g����^sK,}��t����n�H)��K�����e�a-?��0P�|�d�N{ؗ��"fv�X;x'���Ό�9α_��Zv#[8�{�K��l��}�Q5�(����t*�N�#�a>3e��e�ߙ�64;6��K��Ʊﮊy�D?�Y1=��3�4�V df6�0}f�7g�Ydۛ7=<���h���a���w�:�S�B�@��p�l��q���&����*����h�����q����)��������6��(%²V2(r�8.SxЂ��4z?o�Y��p}�`E�Κ�����S����h�^��ͳ��3f:�\��BG{:�U*��{����_9ƍ�b�f�P��
ռ�`�D��ݿC��U����B���K�b�Z~Rq25��7���zF�C/d�sU|y�Iք+PHD@���f&��ۯ_�ꚒEǰ��4�?X�{z&L���1�ì0/�y��T+��;����j�KD@�څ����X
�fz��J�n)�~���=�YhG6!�(�d��]z8kz�x��.s�����.-� y�X��t�L���,���D*ϴ}�x)#4,u��(�TyQ���x��q���7����ǕE���uVNuN�X������Co��- #��#���#? �A��q�eH���Z����Z�P8aέ����2�NAs�_�j�_g;xK_���{��/����/c�ª�ݠ/5;�2X�����tߡ;�|)�N���w�S
oJwD4:�rTfN|�E��5B�WT�<ؙ������X'���ΓE��n�
i��k��#��Æ"zsw]����/�<�s� ����([����f�p�ه&g/�ȇ�A[E1�>w�[8p�}�l���3N-"y�t'߅��_��x�ܨ���M�e�i�����8�E����j��%u<�ͻ_��?���L�k�С���;�J�6/���0^����7�'~s�a��v�~x�O֤�[�GV�e�7g�^�ΛG����MᎰ��Ǆ߬�����U�%����W��o7���Pp��'w'�d�j����o%3���dl��+�3����vr�D'��Q�{��)׎q&��H|�t�7�I�.�dw���RvQmyd�p~���s_Ů���w�s�t�����]s����v�
�=�B�!St��Š��?뙴���z����i�u��d�lNM �-���T:�x��-�yBc󏞚�ޯeT=�VWUUj��?ک�5��3'f����9o�@�!�_v<4���n뜥I��g�5��B<��^l�J���j�gP*�J��^�5�!N	"���u�Ӝ����������z�w�1��e��n�E1|)�U})o�s���qZ�l4شR���d��~�/�0X��,�D�i�u��F�]�Q��F�#�YĜ�%�&�����P��O홟�����t�wt޻�f
�Ea�ofEv������T��%�c���:{���Έ8ģ[����ךª��J��rL�+�N���Z
\ԉ@�F��}��)k;b�t����wz�.�4$?)��<��ɻ����w
o>�jѹ)=&m�1�S4m��~�%@:AD,˫dc�����Zz��-��^f
�I�d�����FX�YS/!H���;eg��Ɨ���Kۃ�~B�P|݌o�2�_�lKCy���s����]��X�Z�W�����C:�t���҃�d0�
�b�.N�=�I��fzk���5��\�B4��r�8s�e,�$^����l;wYTHPtX8�CE���e����,�6n*8}뉟G�tJS�0��]�[1|T��YOu��f`�˗e
="w�e]�w_�B��5�|�v�Ts!����F����">x7��dP���PG��4�6��4+�69�'{M�s9g����݂�a���ԂN����t9-�|S��L&����ҁ��j����3�O��q�����r�)kl������-�]��J,����ٱO�I���{��p�	�$u7X�:���
�W>��m����m�"��Q���ck�a9�V��Y 6Yl�s��=~�b�a�oS}�yƪ�ƌw�Y����NU�0��5�
Pex�S�C�i��G$�����;eş2ݓW�c&���.�6k��I����s�%��z���zs��X�"�Dq�:\��(���a���3�\��0�,�:V��p7�XK�_�<��U���F"��mb�T�tT���>1>�^%*����Z0R-��a�$ �'Zn��ʏ�0c��~����uq����tܤӄ$�n�Ġ#4�oYN��H��.Ȋm!|8`��l����փB���s��'�k�5p�D1=�f����cNn����|^��G�/W�̌��r��Bu�����]'_��DjE�wH��?bg�J�%GǬ-����D#/�]�oq�hֆ��,Hƚ���՞.i���4r *R;�����.�0\�������C��˨ҋ�8�Ӱ���ؓ��3&(�ƣH*q?٦��;K�	-+v���0�~��Ȅ2���=�M�2RlB�k_���cU�mv ���h��x8��w?��"O_��6��!�[�J��Ϻ�*���O%.R}{xZO ��P�Ns�؎6�֦j��+�(����bM`Oy���>ۈ��p�����:}��|{��o�{��s�a՗�e��@���Q8֕�؝-p��%�-��46��yd�� *%��ĝF �r���=�Φp�$� �.���nХTuw$Q�uAa)ɬ�"9B���v#>�a6�ch/�)�б�#4k�nˆ�g;7 gx0��L�P�V �Ca-��G]e���>�Vy�:�p���@kP���~�,9|d8k�v�q��9����]�n���g3xdi{B�k�v�q�<�N��/D�G��߾�ΣP��Z���d�Q��$�s�b��w����@�ԇ�M����IdD�����tjR�aS�߸��>��$Z��e܃�f���e&V�#��$6\3XB����$�|����SWD!?5&f�Tġ�����	~?r�`Z:$��`k��9���h�N�,m�������L[�����1�sJ����xG���+l*�$Ԙ8L4�D4�9�"B�jj�-ְe���H�Ь���h�uL���K���Q���׎&~Ca"-%BWδ����}�շi;V������?�h����5擓G�y2�Ө��zDO�Df���k�o>l�����fs��_��a�v������� ��vRf�u:�oº��������nEJn����;�0��&c}i�{��놞�\�}�'1��������F���DFᱥ��}�"r"!L�N�o�S8����b�Vj,�z��A�+*�
�/�ɳ9��.:��$��Ȣz���G**  ����K;���Byr�ۋ�� �Z�ϕ]c�6�y������N��� $t�wV�=f�Iė�h}[*���\t�2�禙+7�A]Y�5l��M�onZE�#� �G�9'cC�
�j�3��!%`<��`C�dJ�4x�gv��/C���u��)"��/A#%wOZwy٧(�i4�bY��-?!�٪���ic/(���$�vP�N��h���If��i75%@���	0%ċ�z���1,@]�t���E:pk��%:��^w�z|�d\s�X����]8�7���z:� ��2&e�V7q���q��o�;㚱�1�<�@�b�TTۏd��&<���G��4�
����(%�`[�6c]s�}H��ج�̮ϕ9�d_�s _/�)��Z`�ۇg���(�����$/	 �w�5R��4E���J�D����{����3�<�����(��(�/.�2�cU��,U+Ԉ��p�l�%�"̍*�H<�;��o��mhFKF/qƵ[��4;�0���˨��ɞ�Uz��`>ߴ#h �����'݂����0���ml?V�"cd&��d���w9ixeD@ w*sAn���6�Hr��Kf�kJ%ώcHHHp~�8��/"qԗ��I4�To*���=�y�X#�����O���)���ď&���S�f�Pg��LV�3�(��?h%Rm̍��>��f>j���t��:�w������S͂@��:����'���0�e��PM�B�b�D�݈�2�i�����t��M�NW|�l�c)kQ|hBΰj=�s�`��<w�X�C|}�h��̂4�5J߇7J+:,�q�vPp\�o3h��ό���D�rN�jUp��3HT���"X�S�j�����:�;N]��V2D�b��@��>�)�8Zo����D�M�8θ�҉r��2rz��<�ޤQo�⒕�]����kc2��&e�F�0�،g3�A�5nޣC�$8;���ѻ��-u �c��hE7HعW��������n�c��h�����dϣ�̍����nc!�8��S1�O�.���P��ZP�� �X �$1���8�a���Uq;lO]׺�r�[#����DS�Rt��,�7�Q&p���mbU�8{>���İ�r�L�%�A8�S�����{��@�5�e�x z9���B�j��>{s\y� ���
ehYӨ��O+�̳UM�����m@�Ҋғ�ŕx�j�}<j��myHz�o6}�_�YI����O�F���W���'{� ө�M�o:�8��J�LY�[�B�y/8�XU�����%��g!�q�o��3��U��?5��z	܏��R+&���_����~�ű.��o'A����%�����PD۽A�(��`�|��Q"*���+��;�&cq/;�4��P��I�A
�bm3�T"(�'��s���'^X�~�M5n������x��8s��]4_$0���0��r6��?F���D2f��LyXG���凌��	�0��$&8L�2�VM�UF� ȉ��Q�)�.����Wdզ��҅T����"���R��l�Ȩ���b�pw��נ�6��I-��94̴j:��x��'��`�Q��PQM��xCɆ�
��d��-��+��J��4P�>����=s:J���o��ݦ�$K���c�2w~� K�=8`�~޳;6vW��))��U�<�vxdmd!��ϟ��z!�BA�H��&� %�y�� �%�
O]i�'2���>aq��@�h@~[�7��=P���h��83��֏��KF��՗	�a�`�S�xqi�F׹���V5D��)���NI/���vQj��/2X��7��Qz����y��#���X�p��T%���>�
P�i׺m��C�ޖ�t~��m Td�ƴyP����X���,l�����)�T�+m',k#A���::VR|m1ʁ/�77ȶBW^�Ԫ'iO&d�G�H�aA�}�S&�}p�2,�g���԰{���z�Ȩ"��tZQQ�*��[��E(��8�dC�Hܕ���,�[���n�<�eNR�hR�4���ݲ̑�7aОͶ&�4a�󬑺 ��1Q����k}�k�-�����6��ZUI�U~�?�_�7���vGjj�t�'쬹�IɎ!`�'_�VҊ�CH�w0o��M�s��J���i�g������$Exq��k�ϧK�����ά9�Q�0IKN�������K�3%�;p���b�(�E%Y�](��`�)W�O�K�O0Q�s����>@r�0	�ҚC7�3$�Z���e�*�����
�Xj��_Un6�J1�!�^6�Q��%3��Ib��<>bg��W�PmD����@��<��VN�7Z����M�	�"a#��q��q��Y�rm�Q7��$�IB��$� �ի�9SV�J���$�%W�&�¥i靉%��`�A�&$9EfI�@Q���葬�*�;�mJ
�9�_���K�W����`Z3�&��sw���]7�Vj��*]����"�1�	0��������T4�c�����j��x�[¸�\�������̽ H:��VV���$�_>$<
߅�_I�k|���N�T>73e��fw#s��	=a���mg��ӗN�u��.�2��Y��*���Z��KT��]�E�;d}ҿJӜ�L��#�ђ�Tn���|'��r4�`)�ST)O�ϳ��=���aq�;��
R��9�B��$^��W����H-h[�rZ
�s�O>����t�Ǵ�4O_T�^UF\��25�0K��#V�fB� ��'bl��g���]ͷg���_Q������'��Wi�B��fӧ/$*�v?Qz��~��g��z�W�%��J�3����W�꺅��l���W�D XbZ���q�_�y�D�}_��Fr�W��<V'�h0��$�`��5��2�k�UQO����Z걜)�[A��InmiB�A���gmP�-v}��E�>�=ߜh��Ј2�&�DJ��2�Z���o���a}��4a��8�B �x2f���
'��Ka�+���Ԗ|cGɇ���pZ�g8#��U��-����,�۝|����x<��}�c���rY��x^��>Դ��gW�໋��\n�����{�qXdhc]�+�.�3��g{G[0ؓ�.&�})6��[ԫD�ڿ6 ${�G��&$E&9�y���:���۩�?��t]�gz�� u�H���Ģ~F�\L��t���c��ү��z�����c"V�3��v������K%ݹ��y����՛�	nI��Z�̯+�n�~�F��vY�b�_~]kvM��v�?lw��y%Xy�h�$�+�/���}�du��	��˱O��7�	���>E^i �<`��4�o�O�Ǟa�\�/E2�]_�q��.�`�#4�&�~��u۞o��~;��42����ӕ��lNl�6��*�nC��y���|�>]����O�]���G�
C7��\�з���T.C|G|���W���W3�/ë˿�H�_��YtϿ���5�Z�z[-�y�Q�F��c��p\�}����2�(l��[f�O?�*��kzu��(�ԇ%biJf��i����?�欎�sLg�b��r�Hk�4F�*&=�~S���U�fڒ����W��7}*5wK?�$��6�"�x�>7I_���}Â>i��j�H���zm��6����t�����O��9|)�m?�B�u��fٌ�^�Hq=����P��`��Tg/��6�
��Q�:����q�z�O�Kq��%_����:w���m�
�L�L&��<��'f��Zr�#����߸�}�R�Mʃ<�)�Y[љy�f=���E�"�b|������l��Jz.�t�k�m�����F�X�YgR�i�f�_�(;�����/+��j�O��H�:Z�`�i�>����l3'���O�p�r��x1���듺Vľӭ���W.�l��N���<�T_�ebſ�%�Kݪ�ӟ�:?[�����y���q���o4��#��;:�]%�v͙������s�WKN^������{�3i�_�i�G��ŏ��B�+.���C�\ѽ��{��������"U��Q��?����*�0y�jox���mi�s�zi���[(m�q7Ι?�ྜ�/]�����n,'��c&]+���*��w�2�&.�����.p���܀����I����_����@7���܍d�����
� k$ʴ����/ٿ��<�~�ߊ��;�b��q�(�7{����i��*�RP����DJ|�@6�ܮŶ��bui))���S��;��^��p�x�&M�Ih�p�n��.��]�c�����������->��=<�����{�֢0Ԯ����wx�+�_r�9�5�x�>��ޖ�
x�N��HoO�it��4��s����;,�ly�W	�	wa I����r$H�(��.@�р�a %��(��h G�$��9M�����y�}�N��ު:���:@T�*usO�~�ѵ�,�?��*;�*[x �o�� T6�0Pí� ��������;U��ZÜ�[�,��:��׉.��G�C���Do��Q�G�����R��q�tt� x�;�Pb���\F�B�L��s�;� ��]o^����|�d�c�L���g��'L���� 	 ��:o�^�3넞�����yUN	�Yy�� hE���ĺ|}�ɺ�;3H�roqۅ��bA�)c�yt�.-N;�P�U��[G��kfg��r�ׯ~N'ܡ�����
(�q`��K�2�':��=���p'@��+Z�)f9��Cu$�aQ������?9;=lIa��� ����{RӜ�3)���!����ˬ��"��9)֑�}��I�2Ȇf̭Q)��S�e���[�2+g�W�r�����n|/���v������_��x;�[A�����2dnb�<�a*�<G*`���Э|�F��L
���Tj$�)1����S_�����c7қ���aD�f���]�U�면țh�	���r،�
�����@9b�=2~�4D��j�Qvc!^��N��7�-fh�@5��l��.�b�ܺwRA6�獼-����|Cq��V�e���֒����$1� ��h��w�H��)�%�@�^B(4����k����;�7��"��DK�7��Á���*;~�#.�7����������s[�:Ve�Pn��F~�cH�����
>2�H�n 
��|����ϭ�pS�+���:�Jd��;3}�.M�� }�!q� N�6���w�*�;-_x��{Z���1����gЧۍ�i(�cZ��mc�;M���3�o��ꙋWu%a�g'8?֬y�\{~��lJ�Qi��	�(�/�=N�q��J�/�\�����Y�$�{���<O�Y�*�����.A;��Ytz���9�Kq������o'�����A���sO�$�[O�b���m`���?hTO���P/�S��[����[�ͪJA�*?�rP��T�'5���NtD����w����?�L��e�b+�<��V��дqr	&��r#�C0��3��i�6k����6�ͭ���Ke��.\H�jy;Y	��&p�G�}r�JjB��{����I	�������(V2��A��k�n�s�9��V>��M��ʴ���Iھ�Fa�;��	��6�i�Ň�1����5p�����z��ey�\@��M��q-J�y(�F��c���^a7Z���g��\�ŷl�w>z^�vr(�I0d6=->g�P���n�At.dSұ�GW��=�A̒���U�t��v2ׂb�o�0���?M
�mT��r���~�R�>�!��I+������j�ZY.Vw�Z�h`.��JS۹	�����+�s��]��t+痂Ÿ����\���#%39s0W���}����� G� eٌɱS��
6 D�ӽ?��C�F�tlb�.%B�E���jP��a-��
`����v��v��wʤ\r��/+���R؋��.΍5��c���c�|5�5;�6��K�� �{���!`b8�A��	ŗqc�W�!��3���O+��$Y��o�,~j�a��d�	�'��悩�t�nČ�~�Hu\c�;8��79� ��xU͸�&�g�Ip�I�Ӕ�Hv���m���4�Od�����Y&%�D4�U�*�h��h��z��<��c�hDX ��4.z��(��&�9���$���N_?�� �<kg�_�v�u4��h��r����\��u(d�2{�����;�ݭ� %�ƋAs��;��*�L2�~�5�r2���B��S;�}��0��<�yğ5�z�i��%�)Y.�s�Lh�PxN��8.��_�`�A
i�ދ�����X���o߄Mas��������L�[ɠE�wD�"��5��;x%��v�k`.�d��<�F��"q���2�V�S)��}`F��� �}��:�T����e�-��s>�Y|�̷��`=�Y�7.�6�} Ngf���0M��t�w�t0X��&�ϾZ)�"Ϛ/R�R�z:ő&���-1�Á��r�F��[-�o%���+��ߠ�`s4[������7Szۼ6��љU��Q���+�C�D"�N�Z�h������f(18m���:[��?�<�j.� ec����|P�(a�(���J
(��	��tC�3�[���6S��m3+�ZB��	�A�/Ո���*�#U�-:2l�-���g�qb��C�
tR��E�҄僁�ABU|Z│��i�b�D�����m�+ Y���.}RJ�x>����z�����Rb�4DI�F���?��l��:���`��y�6������8�����7��.�iWwق����ގ޸�K|����ދP��f� ��	Ɉg�K	��F�N�����FU�dYQ�q ��0��?�ѐ�q���<��r�CY3�K#v��S�6(�k2��&���:��F����o��s:ڡ�[a����m�;��rPUJ�mZ2�����m*��.�g>�y���9���dV�թ�����F���kxd.𐝯��G��o�V�7���H����z��="m�W���O��Ok�t��1`��Xs�6T{� �[�X�}]��t��F�s-"��DZ[��8i�>��q�nn|�;(�i!�5�r�n|�ج�TX^�6\��]<��(~U��%��c���LR�Y��MU���ٗ��5zv"z��?ƪڃ�� �~����һ\7�i%��'Ui'���m�iH�:�g)�����Y���7�# ������=�U��ϋ͝$\�^���ެx�گ���"�ZQ��bk�>�r�����@��6���!��3�iÊs�X(RRU��^|�"�=���!we�9�v������t.�xk��bk�Q�z�*?���"�Z��¢*|lE|ޓ_���ά��|���_��QJ�yJ�:׭MM��,�в���"��t�� �n��(i���֋j�b�CA��,I���Vy�A��|i�ib-	��KF>;)w.��ֶ�&��H�4?sۛ�$�Ȩ�����~�wP��?�N)���S�Tbŀ*���e�=g�&LISp�CQ 'ը���j�6��~���/[�������X�=���.q̅�$�>�����ԥ��
vw]����0_�+M:�$���x�t�g)-��c���Z\�1m�[ރ\9�
�h����7����Ag��r��mΨ+}�Y�s��J���Ѥ�	��8L�f�5�a�Y@����ǅ;���hc>Ș22-Ͱ�Z�9�b�u+f<��8 �|#��
[��-�{�h�z�ɒ{��o
�Q����`�V����?y�ކC�v�9?��&� ���p��
�i�7	m\�Ǒ<8���#t���<y�`u�I������8�(����Ҵe?���Y�譣,�)q�C�Zc��"��W����Z�A�A�E���a�K:S��CBd���	�Yo��w4�F��8	���|A���#o�wc�ޡ"��� 4���}JQ�������W|�Z�I���`�^/������za��k(��<][U?H�:�5`��K��������C@b�AZ�˰Lǭ�#�?�:+>pNj�?.��������S����-��f�99��aNK������Jb]��@J���y���\ ��[�a�ʣJGA^�Np3�G
oZ�#��/�3�,��XcF}�Tӕ�z
t�u�_O��Om������p�W;�O���Cd;SR8�[�~Y6BW
AZ-����5���iJ�M����h�����[|&.[��}���Ե+)E���{uh���4��MVJq�W,W�l�x=w���/���F�j�E���+�HH�QT�9`un\��{9Zcjm�]W ��ӗ0sQ5�-97�,
 F�k�l\��=U�"&P�'@�_��8郌���2�䐌x�|�6c6���ˁ�����{�KS	qQ�����t��('�T^P0�°S.T��&"h�55>ϡ˴�Ѳ��j��j+�|��P'WQ��.��O97��V��B �W ��_��/rU�G��2���3�,ɝY������
��)�bNtf�m���\�b��;Ԭ�IU q 4�di��񦣮�����Pv����EF�Y���ncb���څ�=]��0��]������FTN&���>�+�c��7r�TӾc�R�I÷�⛔o��͡�w��0��56��Mb[��i�o��,�$�3kȟY�^��[D뙔��=��ː֩�<�)6*���q��7�f7㮕��X�NxZ�}��������I��[S��+<3�z���La�x��&�wy촻�V�K|�!)����A�A�FQп�}�u	���V�y&��� AbS�y`���$���z� �P{����ܛ�O�C`�G�IW^Ć����C�E����V
�Ӻa��$�&���Ȳ�~%� z@,������(��G�z�I�S[Y&��.w�7�$���~�jY�=���t��h �EP|�g�6�5
C�#�B�g۾?12}����K �*b��9�����]:�ty��"��{�W�l�\b.�l��Z/�Y5��Ż"jf.w�����C'���靕h���)��蝄�Ût�+�z�D;�(��˛�j�X���Ȝ���c���
��|Q�t.�/���]����9
��I��lX$p#��l��:�f���*ķ�0���\�ֶ1����xT���c�t��(����Ǒ�_6����JUwz"U�g�ޞ"�r<B:*���b�Ý~�7V�)]U����ƏF��#X�b&&-`Z�Š�����克�p�2[���j�����`�LrMԲ��+/O6'���t�.9�A�] ����2Uv>���n;���XI�h[E�_7<��	���$̣T~	PF��"�Pv�� @�C#���-��l�A>�`m4b|��I��T�ZBKH���E��<s�pʷ�+�uLfg
�hz}�G�5C1�Cn��9?���N�m���$�n���ST<�̍j�!ΗsR�����H�t� ��Xnsb�{��BPyԾ��le�;�0H���p�g�T���>te �.TauδxFR��gq��X��b|N���**e捊����E�b��4F]:Ɨ7�tk�Q����r>��Ƕ�'B� %:��_M�Y,=���+�yWE�j�m5��<B(��K{��	u�2���Cb�<�QJ`�M  l��e����x��.��m���K)��˭a�F���}ݵ?�}g߽������'��ӊ�K�f����/�"�A��V�����ZϬ|��y3�T9�;Q[WY�v��V[P��Q�9}�?��tc-���I�jhlUFWڱ�|��GWP �turZ�b�+@e�����#�tn%��Q0�H$�#W�n��O�MhBH@��a�]"�ߒ���L2��㝏2�އ�VqS��1�EaŘ�SA�][�Fy�|$����B�h�Y�a��� �qk�q�ڣV�w���g�@�s�ܪ��3�N�~��4�	�k`e&�j���y�%P��
�r�e��u	����%�ǩM'T���ŌV���xz�ʅ5�L�*��ހ�tCVG�t3O��N��ZOb1Te�k5&�3����G���of��`<i �-.�9�mk�B�r ����
�U$��?8��ip�"���N��R�*V�ھ5�k���wS6>�-�k����3Qk\s4Y�/�a[W��1z��M�
w�.�{[��>�<�L���9��Z�G>{�������̇�&��Ε��߅� $��Kj6z��x�LT�,vd�nG��T�弾�-���O�k��.�n}PA�-Y��{;�V
�[xԡЎj�ۿ�(�݊ �]^���Ox�Z�44#�ё��Trb%̟�ڣ���?�k��k�+���T�;���F/	-���o�kY)w�z[^Q��HS|o����|E=j � �2(Ot�la�X�*�Q�K�!*�+���ՊX	pʢ
_ N^�9$=1O�`��l����tZ�U(Z���a��)�<}��z�ud�34FK�f�Ǜ�:��͍�`��x:B1w��Mq�K�mm����V ���<�2�?%����\�����<Z���#��'%�A��5P�o������/�BW���p���9����c)��A���咼D��皩Ϗ:ax�F����2_����3��I4�yi�rP��OpblW��/�p�|�(E��1�`�S�Nv'�g�EZ)��j2޼
�%@��sR�*��6�j��)t�A�h���;��f� Qy�N��z�i<'ds$���8������p4�hi܉ M��[RC���(�!�G��<��zƢ+m.�×�MN3�������z��Z�:��)/�GL8׺��\��{��m_j��c
�]3�S�}M@#��M�oޙn����~5AO�Qs����[j54eՕ#��+M�x���Dᕝz�|(�����Ö籧��
����}�����
j_.�_����WS�b��6ɵ���g��Q�E��΂MT	�]z`�@�>���F��#L&��BBg�V�P�׀TF-ע�/ݶ^xE���&j���~�����z"Tw������ m�x,��<���agN}k'�s~I�kc����2tŭ$���<,@�^4X��gsm��ڴ���6ir2Ci(�cy�]Y=���4,59M�s!M&�u�j��į�"e�˒��E�s�y3z��[g����JW�f�<�$Ԋ�P�O"����i �g�����d7�=G@�3�S��8-*��nQ㓔��j���H.���E�'cs�a�1��z�	%��:N�@7|����S���qP)2"N	۰��'���T+���D��P�W������j�!���V�#m��P��.i���Y����)����]�e����2'/�2QX���uTr�^�B_���l���|CGZ�o���(���9�t��4ڌ��KkA�0�\:��J�5�[����(�2�R��g�����k��we)OH̉Z�eT5n�V����\���܀����&�5�`y ����k�� ���/uG�l_�$޿ڙt؄}#tk��3�JFX�/�������Hxx83���&��,��9�"@c��đ�#�QCPT@��ϋO
���[@S�����g��r�
�:M���_Vv�* �q-U�hk��U���}U�����:�*����'��JrkG�),����p���OPHXC�� ��?��?�&>d<+}Ғ��,�r�}N����������$hz(��d�8�a��p9����3;4j{�l�N؄N�� "��[���n�6`�nV�����uq�k�����I�j�ZOc^Г+z�y�=w�خ�63/>�DN~@*���0��
�b>�:��i����/#o�yJ�ƻ���X�R
s�)�}a��Wl�?o��ZF��7=��E����T���
��!���ܾ̩���;~��<Q Ϭ�������B���cdq3f#_��yt�q-�A�3�[�� &�@,���Е��釾���<+�4�0F��ǤrZ׉'j{�|�6˖Nz3��;Y�ؤ�6���~�x�*<+1�>kW}�x���� ��;��* �QZ��!�
�ퟎAVg�}?�_�3}��}�o�k,k�����:���<�6�|y���^�D�G���i!zWv:����}Igޥ��޻��߻Ln�;V%�AW6M�=P�T��e1o�r�t�H�0���F˩��8�ƞ���}e���l�es`�����N4~"��~D3�p����i�r����Wֻe I;ɛ#�?�3h���`��B�<��xG靾�Y��i��S���t������������Ç��#��on\۸=ul�
���V�^yn�Υ��N�E�<�jN(}�����Z��|#�Iۉ��G�d�`P�|ƣKf��&&��m,E9 ���q�s�i�OB���})�f����ܓ�Y��¦~� �L���=kZdk��I̾E"p)�G&Eg�/u�Dr�r��o�2~�$���k�SY�,�X?��s<�����T�:�S9����~hzϖ��/t�2T�0��H0)�r<`���BT7���΄-J~h/���|Z��)X:��)� F~s��Q?� �j�E��pg�>\V������f�$�-"�AWj��ܒg{�5:!�굺CS����@�k�B{}���ͧ��uh]Do����;��	���[�k��꺱����,3O�U�y���Qh��p�"��bOvl@4��U�����^+MܾS���`8��L�NeI��D�&~!�ɺ"�_05��GcC���/�L��&J�~�����-?�S�o>���8|��] ������k+N��w0�׷�g��j�f�90(�:�0��T�Iқ�}:�lP���B4�_�wh�g�����Xv��� �Sw�8P���ߴ���}�����H�L�\)�O�Õ%���?��-�,���LH����ɥ��?h>��KxWc=���-����|�h�����c�z��X��W'�C��G\�!)kwFg4ɻ-є�,��-KQ�o��$�ۺd����{�`�όv����ȃ(1h��ӿ�"(&�7$����YH��=	�&�Z�k{Km=�ki�A�I�nY�y'gﲵ��P�.Y:�r�(C73�2V�(��Y��6Ֆ���M�) @BC�l�fySO����R��L�
w\�P�x���j>�ܫ�� �Su��*�/��ˡ�|�ȧx:��_�v��������g �}?��$*̽���df�&�p�fk���1.���ߡ��g���e.��-�'�F�e��xa�U G�&��{��e�Y��#O�F�����+?��l�x�ч�P|�O[~iWmj�d1�X
����:d��Y�W��#0�����u��}��������j�xZZ���a��LL���x�����/o�5� �N��sa#��濥} ���b;iM��2Y|�j�h9��ՠ�;�v7����9���F�ŋ�FP�ňM�"�X`��J�v��eh���E���2N��oޞ���|���l5�s�e̾�9�N�>~l����{�Sq��ktT�ڲ]�O�_�-uXw@Eҝ�n{'�
�;A�����sE�V
�ei0i��*��1䶢�cxM����E�x�* q���l"��Sϒ6�!�v~�d�\kҗ��F�Y@;L�.�����\"k獊�����o͕@�����]aVi��Ȱ%}P�:��v��#s�ҵ���%�{So;D�I:���W�b�M�
�@��� o� (��STF�s�#U/㺸g�6��n�B�}>a�����tF�Ү���"law6��Z���q �t�m���D0C�^�� �	��Լc= VF�D'c���?:b�ݓ�FU���8}H �;A'�	c��1|t 5VȔ�d��:�j� MTj�u*�qu��V�z�5sU%Ū�>�f�`����-g��\1T�F��K����{Yk˦E3y���@��V�V^XE�̓xw��ؠo����qH�"�����1�X#��Bȕ���?'��,%'&�,�e�S �MN��S�5�B2��Y$[��ϱ����������fpʿ��v�~��� ����h2UV���z��UQ�u#Y�k5��4yи �U�վ�8�R|U1� R�իrn�3v��qq��#���Q)+<�P�O�Ԡl@��׊��$X����}�
�*�X�J�+��;7�!�W��r����|��?wd�:��XB���X=� �Y��׵��EUW�NQ���\TX{`���ʺ��3*���v��j-_�Y�^���՘�|���e�<=�$�x��F�O7�͎'��:}�kE� �Ӭ�J�_�+�G����>���@�V;��� ��	e�k���PD��}�{�`K�%Co���N�=�YZ���E/��PJ���3�S���D�DF*|� �ל�u�����At������pb�u�T�s Fݲ�T���躴t�z��R�P���o:�����`�i�Ykؓ�S���x�L�����Z�2�f7J+��i�#S䷎�&��ǃ{ZP�L� ��$=��S���J�wc��{,�N�D]I����n�p��Ϋ���m<Vf��/^4��C<$�NR����i2b��J�� ��[J*��l�@���@�S����f)�ߒ�H.T��j: �f۾:�g���U�|e����:��瞾���e�%���ST��ݞ>�ڝ��?���y�ם��;a��������_�P3]?4T �8����OvC��R%�yr����U���x*�<�������!�,����m�,ѓ����d�[��.k5��J�/$�]��Ld|Ʋ���F! #	�����.�rφ��"�ӕsd㻟�j�k�N��tg�j�=M{�kS�޻���"�R��.�;'F�Ā�t�1VUKƥe��k�� `��W���0i��b$�nYZ��_���{ s�=�Ǿ�E�d�/�4��V=� �35��Rx����e�EȈ��(ŗަJS?f����~������_� .̛\�j���#d�t=�t@"���dO|TC�T]�b�"Kg�5��ŏ{4c�p���mb�;0Y�n҇v��JS+5�Ӽ�>k	���@���V)�� Y�c�'�Fl�I�S��07��1;�!#���~�'����FxB2�~��|~�����/�#	o��н@ad;�7K���?$��3�������;ܾ۠ ����a̾�F��P6�}�v�&
�7�mZ^ϻ�I��H�'!�3��S�O����gR`���E�9�?�A�"4�O��Gn������2LGC�5�n� ����fw���2�Q��"r.����Y�x��rVCr��(v1��&��H3°'�~�-�g;r��8�_ȕ���ڸ�Y�G�����bc�ul6S��l�:�h���~b���Ъ� )_v,��s4�S�� ���(G[IP%�|R�H��W���C+��f �Z��݋}t��!P���ꇹ�����x��@�˚�d{��z>�Ĵ����T�9�VL�Xp��+3�~����L�F����0�~l�G���� $��:��5��[�ڙ��%��>�1�ꜯ\x�hp�8u�F���R�1��͘�Ud�r
����𤃊R��s��ks0��%�6���p�L����d��CNU$��ڙiT�P������)�k�ݫ�ɖg'��8
	9��Sm�3�Ͻ&�+h�rL~�T�W�M���/�c�A12�%�!�U�s~��Nߢ�u,��"�>�Ƅ�h��ߖ۔�I`�؀��[�q�����Dm�r,��g�� @��W]*+�s;�����/�9ܲ��qI��k?{���A('I��u�_~[>�n��jP�}d��KP�62����8I�'Ȓņ�lɛ���y�AH�;ߜ1������F9��N�\������P���^7�}��-�p����4�jD�zM�A��A���|��c��d��U�C2c�4�CU3�y˵���.I��Ԇ	aJys��~�ct�F�R%�]&����)���Zo�5Kn�������L��z���3���מ�'�M\_&�.z\��)��%siÕNUc�d#�yS�Ut/E �ۗ�k�d�%��@4��X�i=��$�x��8E�*�$�ק���T�춄r*H&�v���l�&�?���Y���?��ťC��7�:Y�W�b��S�=��7�AO
�z�ZMƋj�����wܝE��1ݤӏ���\�ƾ�'GEJ���^��?�2���c`{P��ŧk�mh\�*�����1���ϛϜp-��_/���a�e�{7�5dc:dF
��&JiL�>�+<F`�|�F�;^�5Ӱ�a�!m����0�%h]�B9�Y|��w�TY2�27����"���Vf;���,��ǡ�f0��luhۍ�kXǀ�j&_��CC������g���E���$�8��KM��;6E��Ӏg�C��p1Z!�l��]���4�~.@����~�4�	�%�3}�h��aas���Ճq�u�x�U�6�N5q)��������,'N�rAG�=3�}K�ouQ���ں�0������n�v��+��h(8�+3�i�cjv�_��mȭ���LhL�6}��Nl��me��A�H������
Ŧ�]��­2ܪ��3Aˆ^�%����n<��F
�6w��F9�;Ц�����!�z����x�t�:�=G&>�,N������o�L��w�%��OAx��S�+�/��a���x	^7��t(W�k�_N`[<{���.w�ѥ��0�'�kᆬ�>Կ�'��z1�g��C= Pc��s��^���6GT�C���緖�۶&�v2�-%T6��y{A#^p���� �.��GU3�=��z��%l�Y�6[�h�f|�}׌i�B�^q�����,}�yB��G�mi�D��"����3\��><.�(-

)}mkn�]WD+��;6v�C�=�C���G�t:��& �ڝQ�`�����bgP)�_$.�n�-�;�ۗ�?��g�`g-�ץ���չ�\�{�Yit�a�Rn\ PX��9v�M��W.p`��-�2��C��a|m����2�*8P��,��N��s5�Y�Y��4��G헻 	OgI�T�#8�d��,`>mhY��; ���$�#����.��*���i��f�5������kT]k>JV�h��3���	 S��Y�{^�
��}��:tsm��ͤ8�0=f?C���n�L
0BǢ:Ty�b]:�X�0���CxZ��>{��%�vvܧ�s SŞs����)�!���y-�x�Uq���C�}O+s�':�t��w8J?��.�*.��Fu=tMM�r�yC�p�*С��"�(�B)O�{�b�߇o9�]�6z�]�� �N ������OA)��:9��e̺�"6a#@���^U��&ɛ7����=���,mk	HU	�u|�H-'��'uac?�D6(My�2�v�����<4.'8��, �Qm�u�h�� 8<u&�r1�_��������Y���U�農X͢�����=��A��z��6��<n����f 	p�� ��L��N��D	������i]48�C�]eh?�]_�uTi�X�����_�wE�j�}tm˜=���&�-�o7�`�AOE�T��k����h�	�~�}���`AO�h�꺁��S�f�֒ �����݄>tI%j���s�i[�Y�铷q	�%�U#��������.����ã��[W��l���@�
��t|B#�L���w���,���"\��]�?e�*'��޾�.����x>���p��]'6�3�#�z�
iA�;�Gχ;0�4��t@��|�]{zs1Vg)z���xق�X4G%�(��B\�#��q32g�C��Aͻy5���m#��BL��4t��?j*�%�	w`^d=F�XY�����m>�� �4ӊԸ�؆Ǐk{$����D�����Ro�NS��:RO]ݫt�����@5��h��)2��  ���jv3�������]�U#�k[�x� ��.za�E��ѣ�q�T3�A��^%�*(�;���vD�o��X�eI�ɪ� �tWQl����Zw�R�Py�%hQ�Ovs�ݠA>�K�P=�{�+{��Ɔ���۲���$ ��9���A�Ჷ�����	z�pdH�v�C����OǯD��=����Z��� >�\"\��0�X��"d2��*=�򫸂��ZM��2��^.�������TR� xI�ŗT����T���>���	��~����)�|��Ho9�4v�WW������T���(��z�\�����K��{�B �V�����.�j��B����JM	��<D9{���ă�b���Ϋ�?�s�7@��f;3&�OW�8�uJE	�Ԣ���ro�a��J��h��+�a-���o9e,\VOu�^�"�Ǿ��1��,�VW���ۃ���8�U����7��_�k�qޭq�ؘ�w�2�jzxh �v9�9��dǚ"[M�[�<0p�^��^w�������?��v�`�9R�?Z��Z��bC4��+���������S�F������K�9�cɀff^+"]��Ž5	���D3���c������¸L�u�/��E��!M�W���W	��_w�{�ǔ1$:�� ���k_x��v�4�8�v�ȅh9�n���������m]�z���Ɠ�ڋ��-ZI��L���T����L�1�1sk�W&�U������+��G+�q����1�B�N�ӵ�H�˜��Xt	�.@�]�4�2<J��Ƈ�l���U ��o�l{�?t��o�aW������?"��;Q1�Yx���� �$�FM�E�1:��
��S�� >�D��t�E{/~���.I'�C����j���'������\��]�"��!�A�V�M���[Um��5@$��u[a�1�j����e^-�,4!��1N#<���\C	���.���|]���fC�I^0���.��}���/g䪱%.U��Q�p��v���V.�:��:��J,ݣEn��6��}/5 uN�7rW�.�"��z��M�����ޅ|f�>XJ]��2�s���c�Cpo��2��6����>I���>�|�;�#zR���X�K����'$������1�B��$ŵ�&��3t��(�K�8S���q�������ޅ�ܕ��c�T��8B?̾Y��y�{���f|�,z}��8��M�"��Eq�>ݞ��z�~�gh�v���ͼ-tF�ZD�t�n
�g�$��U���c���Gy�l�zӢ�`��t�w7:�r{k ��8��W��>�s2����9h����%���M�ъ��F_��m$L��-�e˳�����z)��H��Q\A\��,�g?ǜ�7�i��s�(�etܒ�5�����)���l��F�DC5�{}��������1,�J��2���RG)j݌+x�F�0C�8;�)��+xn��p��(�Y��*��3x��,�]��A�'흝����O���(s��¿OV�W|�x�&��A.��ˡ��v?�1	7��s���'Q	wc=��LN��_���B�}�r�g�2Sz"a��͠��<�3Q�4[E�d3�hk��osO��Ϋ�A��ߓyQ1sx��~)z�������w�Y��ȧ���H���?tt�/@�(�@�oekH��N�`�4�4��
�Y
��;(g�O�Sy���j�����ST�!h���\	��H��gv�C���/��ǧL��#\A<	 ��Q9��%�d1�7 �%�wJyz��`�E|�o�� h����,��C�?1{Pb��
i�d��po�~���p; �s~��z�]\W� �]��owe�bmf��j��H��u�tu��X�ZҶ�Ƥ�Y0�Nj �]/T��}���`(G���C�_L�Ŀ�A���}B�T�]�Ʌ+Pl��lx��$��L�`�.fS1�^.��Ό�?�̍ρG\�^L��K==o4+(��W�`�]e�?��� � �'���\n=Xu��WO�M����(��`B��ms�!a�����a���GU�d]H�?�xk������7޹�o�6Mt���h��W��Z�e�/�7���v��&�n�&�£;4�sR�� �� �Z�Z4�:3�{��I������i�p"���c�# Z��W���9��P��D	�Z5�>)�1j�R�o��_�mi�>V�T�IJO�����o;���_�8��9�*�;�J���?��#�I�Yx�|ޠ��aqU�e�Qv���Zq �����0�Uz<�a2�j7��R��*~V�.��@�se�|J�5*����}*|��x�����'�R����ePs��̌���ypPo2����uj47+�#� �Ճ.'oG����~E���K����x{���(�L�9y��3 �ܾ��e���g��+>��l��m�[��U�����/bf��R���P�yI��1v�򵰏V�/1�v�slDB8�C��:�j�]*Ǜ�q�pK'z�҇�r�k��䵇�}ȟc)W��;��i缍[�l1�NG0��K��LF�[��pxi8���eEK;[���� �Jq{}�j�Ja����Ըt/&/�);��[	��-7��烓��@�G�G��j��`@�J�z'$M*d��YBW���߉���*���a�'�D��_�k���D'�h����ݨ;�����b�2�РNWp��,5�o�1՛}B({Ӿ��l����D��e�ш<|
�V�8@=yfk��$�'�S��
'�Y��WJ��s��P���jo���*��i��@r:�Ќ��O�<��t��� w��8vQ�X�4�� @�N���1�ZG�T���#��j���p-#O�[�q�I�3$�*�D�KuS��;qU�%��6�	 Vh�������U�.�R�`Kv��ҵ�#��^>#]:W�F�E�������b���0���x�Zw�oǋ�Wh�ӻhx����o F�s��H�����,��"�=ZwKR��C�\v%��� Y"8��-����M�E�ȾN6��E�T�2�I--�Dm�"s�*soЩYe������#�, �����Y������諫�ρ�-�Z�|�2�26*[X��5Y���@R�5�v֝��0���vj�h��eZAL��T�5�NRsZ����U�����1���%@��ꐹIe^Vr�+}W@�G�nV	.�NbwV]Ѭ�'e�=��  �$:���5~��7�LŬ��1"f ��y���h][;��w`G�>�� ��v�x�Y�d@�8r�H!��7��`}'��5s�g�;�q?��l�)��h���׊����7��W��ʷ�J��
�n%�1/�o��1q��[�����]W��v��M�{��O�ς`t�P�3����?�����tGP���'��rxz��o㥝���bx����x��|Q��M3y�� ��>��� o�?i?����C������ �^f�m��N�*�H6�_�0����,��2�H�-M��J�~A�\�M#�6z�!����,��?�ॹ�0�m0(@�Ö���{҆�E��2�k� a ׯE�0�����oA7����1��P)�&�&/vڰR���@�4L.���pW��+o��Q�	�=��Qu2�C�8������ȩ����l	�߇�u���O��+^�#.~b���	�80�����k����Q�w!���ʵ��PC�{(<r�e�5i����w��澋��f����#B�WA�����/��4�ek�&E�rzJv}�8n2��>��m���ڣ�.e�%^����BQ:�Ig5j�Hm�Y.קdz��ރ���%F��l�E|���3x/:?���?�A��L<�k1�)�_����C�!%�Ex;�L]��>{�z��V��k<L�~L��2$6JdӲ�	F�^�\|BrJ�p��M��[]`˴G�bA���U�"�M�Buq�N)�SO!� ���!�)�x�a5�x�̎_C�#�q���?�� �P{�YV�6o����!�s�t��RH��0\i8�;��u+ȕ�=(K�zyGM���9Rf�$=��I@�rm�ZԺTLJu�!~LWɶ�ӄ:F���!ɋ��C<����)P�������MȌ�	�U���A�@�N�����NlaBl�9�*7�k�Ϛ����.�k�^��׀��>D�x�I2_d7��lr�#�(M��m-���թ���ܓ}�z8�Q�@7bl4�5Fu�kQU�];ݟ=��0�H��b{��N"g���!{|���'*{Q�T�A<��J!Df Ou1�p�����;.��`m4߯�sy����{�B�PZ�Kl��d�]R�g�F\�T��y��I������@	�ѯ�����%���
g��;�g�:-G*�͸�t��&���� ����~l[~"���XN�pDHW6�M��x��?S(R�*��
��|��<��G��I���(��^��1��R���X�x@��W0�l~����+���w ��d?vɕ�j�R_8R���"���ú�������D,�0�$��	�,a�0D��T�nH�֖Ѹ�LQ��"�we�����)�Q	�lql�����BIr*zك��5�`3�( ���-"�z�/�1���L�7^d��O��&��B��j���p���FV��Ld� qP�k+��@Ԉ�Hę�������.�`�`&'�|�] HL/��h�cL
�ꈊ�+�AX��A=�'Z�`
N�9�����$��Iz0Vg(+V5�;ޏ]_�#��k���X�H X��8�ߑ�����Ü5n��i榞�ѐ��Iju��_��=X�EĀ�O��S+S�;��IȹX�H0�����~�J����.+��t�Px-���-�����n�z�ɔ��TJ�sl(�\�8�?/�\��ᶝ A!�Ny�� �q�Q�K�G�Y�XNOW_�kA9Y�^��^�g"��3��ް�uw�-K��w;���*m���C�ͩ���[oԄ�A�����|�Aj9)=yN&O�^��+��it:�8y��4�lM�|��uB��>���'/b�%@2���ς�~�����K��G�����/��v�R���~�e����3�^#.\Q�"=r�c>Y�2(������L�)�RZP��ӁY 5��]�QS�:�Ƞ�9��H��;�����K����P��iXF���ݍK��	�QY?���2���h�i��&.6�K<6?ę�R]9v� �!#X`e�鄘Y�-��"m����.�_��E��L]y T��Wn����M����J!B�� �}Ϛ}���e�ʒ*�ؗc0�dg$�m�[���{�,���ߙ�<���<�{�{R�Y�W�'�e`��_3ƨ2T�#��{Y�A�8G�8�(ѥW�}S>�<	?oJ���K��g������kod���}��'/g���O�.�"@������9V[�5`��M���2 �̄�e�\��Xߑn��r�O�n�o��R}�}4��n�g&+*j�3�\m\� .Ȋ�;x�P�'�M�������F=��*P���Y�)�L((�	�� ;!�l�b�+�W 4v9����1���;M��f:=74�XNw*�{X��?uC�U��$�GrobH]C1�Gw~Gf=��h�!�G�(>�n�>}�J#&4�2�o��v��,]�8d�S�?L�r\��gCլ�_�����S��:��h׋��	��e����v��S@V��C�}�������o-�U�W%�'T����v�юO�UĬ��_��E)��ۻG,^���g�w��6�y�	PL���6le_��R������"�w�)s�'i��kb��a��﬉��`���f�c��0������
�
qHD��Gt�M��.�k����3w�{�3�:��K1��.�2�ك�:B��z`�m�rS�(@:�0+����W�lI����n� ��>��u�S����5�t�k˟g��eÚo�]�,��ה7,�o�����zA:�(.<h�3��墣�E�_�>�������g��]�ډ[ty��_#S����my.�& i=` kh�\ս���BnۦO ]8	�IF<qg��还<-��VS8]c	����?�^����	0�� q2 $ׄ����Nx�ó~�Sp�O�9q�����h�_<gW�|�Bp{��%tbn�N�ȡ[�]�@Г����&'�u��D����������f�Dz;���O��<d6���~��1��T`��ob%���h�S�f�*��Y��̀@l��qn}	�?����?�t��'���1�n a�7����+o�N<�M��1苒!`���V-��o��՛o�T��캫8b!�n��6=���?V��0�*P	\c j��*���g�\5X�V|l0S��$��]:߹`E�������E}I�R�(4(������[��-c�y���"(�X҅�����E^î(�ѻK��+��_��������Lx��~�rk��N�0�䭁��;��6�_�/�< ^Ȗ��:|yK���Y��`Axp��&�?ua��4�pJQ�����	��@�p˺z-s�?-/���egt]�}�+��wf��Y�Mp!vg�/�jj�J6�15	1zg�����-�ٽ�<	b�?i�4�5^���U����`<�fy|��mP��U���6�0�	n׫Q�x��a�����1A����A
�H���B<Th'e�ډ;�t�?��GН/	ӿA;_sh����݇�;?}�[4��{'��k�1:z��
�"e�7�m���@D3�T���{�H�`
k
^՝� �'y�4<rwpu~Յ�`2{ uee���hg��|t�\�t����2�C�Ԑt�b
��^�D	�!y�.��p�{
��.g�R�cU�-������ۑ�y�#?�KM�Z2�駘��Z@J)V�\��=�{0(�ï�*�������Q���z�t���|�.?��ea]��p(�	�3[��:�Hh���	�[��(	�~�^�ⅴ��������Lg�H�6�a��kW��Ar5�-Y��L��y���FPp���f�nhɱ����T�Z��o��~^-!��Z�S��`UP�ϭ9�֡���K�&�������1���@xѮm1�n?�s����h;��� �J.�ܖ�O�l �z�5Y�8�u������0�?��Z�etN���i$�\�	�Nm����6�8x׉�BM�w�JѰ1`0�KW�:H4�Nlm7W~E{70�}O����0��	!in-�O��;�)	o��J�f�LR}z	/����4ޣ����(Eð6`'��E�0�S�㒥�]k��.��<�+_�$2�Mg����A��:K�+�x�@��G���q��-�'���%z:�t�(�>@ eiZ��nd���|j�8��z_g�/�i+Cr����4�(���<�&�3� �p!��kp>t]�P��#Q�
@Iç&�,k��p�T=�cP�=H*Y�$���P!�����U$s~�5e1e�Q&���Y���͙4����럿<��x���s5��O����G}9��{�����''�+����>����W��Y;'�&�8?��B��mɈ1��|7�P�p�_"C�6;���_{{��w����:N+Z���>L�?>�q�j�e=���a�z̴p�|�|�~��1>�g���>�xtr��	tu�S��?����:�P�k�|��l�c9�kS��I�;��dA-�n�>=i�=od��z�,�͖�1�j���\��8U�s��>��p��^�Ì!��:��|&t�LV�!\���ӴP�8��q�L��7,l4{���S��p9W4=k�WR7F����: t���Um�8y�뾧���0-߫u�9�jb�㏤®�M�A!)�"�i}���ۏ��x�&�i�38G�q㫨:�
�|�Ęf��q���О�*��AT��I�!��Όxbg٧~�l\ �|6{�@>!c{jpJ�U`=o7ae�'~��PPdx��@���� ��oo���L�
�D;����D5gٱ3��A�ί'�z�J} �FL{�9�)#cB�-i���E��AY��O��W�����������gB�s�mm88���a.�f̺��1<\_L����5���y�Q�������1�tl�9�q��� �%�:}f:��3(F�*.��i����;�Omr��M���LI-�� l�	���v_�C�N�u��B��0l�����O-��U��Ni�֛I�嚴#��c���>f�u��E^�>?��J��ar��o��"�QS'��Qm,�~��?c��D�~SU�C�eO��\1��Iiȟ��䞏�M=rVrȮ #q���������ͦ�M^���M�F���_gb��Ͼ��Tj�p��+��_�{@l���Gڥn��e;<�W͘O�����4��z"?�C��P�cU����ZgĜ/�����[�^�V�˶<[�X�<7T����Q���:�|��d��i	��Z�î�#��}f��=��9n��������{Fz�9Jg�����	�U�h���W��N��d�T_�x��jd&�̨-W����Ji�3i�%g��9�1�����6e<����t[I���,σ�n�釅@tY�co�˗���)�YL����yǢ�5i��Bx��@|+����'+ +#�̕�Yd7Z�*�Hg��L�د3+Ε��AH-�*��C9C_�t�cj�UB��'����1�=�% %�� �^��퐳\�_����M�}����T�]���+�"V��ES�$'���;*fB8���	�7|��:~M-V�������VN��O�!#+l��2�f�������:�a���,,r&{~a��b��gw��ȉ՞�z���z���@������%O�N� ��}�/�	D�! �M�d�/��~eǙ�Z�q�i�3�?�Ƕ�ݼ����V��U����@b��(�W�w/�/{�o"t���=�IQ���*8��+�
�-���#5$���oVlu3����U�����h��ح~�������gߊ�iٗq��ᩯ�5��jo|��4Y�}�e���L�t���M`�/�UѼ��N�<	f	��!�1 Fq�I���IK����:VXY��~u�v+?�&����V�.�נ��l
F=��i�5"M��/b� \)�+����S{�n�O���k�~�bZ&Y�����x]�o���۫?����Tbh��`�kZ*�@���4б���"��}�X��U��Y(���a�K�vU��8����X~��ɡ�:|�2�AV:�.�)�KJ�����+��QǘX��j��ט��B0�v�%ݔX����zI�����1�>I�*v��N:�T�S�>��}Fc��~�G�d��Q�U�,�m�O�,\ɯ}A>�My�r	4X��M�|��}�.~������䳎�UA\�/�>ԑ��w�v\��3$�֥%�3�Fa�%��tII�2��a�b��6���,�=?㱬r�-"22�#%�����m�.4�_�2���|e"����\_@/��������C�d��C���ȴ$�۵��{�8���Z��dx>����9����ۼ�;��2ۖb��HǬg����Mj��#���(lE�^pm_6��шL*�(40�W�ǯ�=�/�"K^����?Ȏ�Q}�i�rQ���r�Ja��pJ(E(�O�èˤ���?j��tɻ*1�3CQ�ǙV�f�Xe�7����4X�M��zm��N�;1A$��X��=�L����h$^'hB�j
 A���+%I�X��£}D/dl�,�j[tPRHB�N��u�9�l�����1����4�_����ev�o�D���P$�PXL���ZiJQL����Tr|�;���1Ӫ�e.�-�d��7�S�6�Tj�s#u`�a^Y	��o��va��<�5�~��Г�	�L�E�\�a�W�D���ݶ�M�g��P\c�,-�أX�ƚ)��`��!/\#���wC��Ċ ����eb=��<*�-cp
td�u?ɕvO�N���v�1�jgEmyE(���\��a��G�Ω_�Hˇ�v�
�X
n9�hj9�I��5Q�z�l��5���>�j��A}Q�0�j+�O��PjȆ����Ga�����#֑��s�5��$�7}C�"b&�Ol��'
�DՏC1�� �j��C�l�uGd��{����8x� ��z6	��nTc�ρ qr�k��ZJ�5X��A%�=)���}����ȩ� p�c�rn[�v�8n�j^�@���`^Y�3pxe}��ez�1����Bmi�֛q6���)�я�g���G�+j�}!���aixW 1�Vj��m��z��Ї���,)i�1��k�JdW�
;&��m�Ѯ�l_6KE���yX��x�v�����2�p�\�A潸��P�\˩��G}ɳ�Qli��m'��p�E��хGNj��f��e�j���1�fim�� �T8��O�E����˿�6П���B��q�='��������
!Q7E�4h�b��e�Qf�Sb��D	�� �J�m�hj�Ciq�����\�t�3���6��H�l�� V�c�m�DK���:�]�i>G�L��^��_Cy����v�L.�L~t�K��Ӈ�g�t�C2��!g��sdK�*j=3/�*1;L��<��=:�|��)m���4@�����"W\'h����-���{���c�y.�9��d��緋wTeM^H��Ik�m"{�����ph=Ym��ǩ~���yD���L#9Z[}�z�����y�W&CE��u�O����-�.�pð�/�N���HG��N�~�$r������%2 ��0o����C�B�|+ef���8��L�J ��7Yq���t��om^6�K}�>wO�X�jq�_(�z�X<�@"�C|5��d*�rl�E��[��ֵ����$���:C3��X�z�F��d�<Gy^'���L���
]]3Ɨ`1��GTo���2���w�e�hY�>/��^&����CGHA��1��&��9�.�e���B?mZ�cnS�����P��,ʮx�Gm�yMh���%��n�d�Q�,����/��h<q�ʹ�+nbO������1�L��e�-��|<4��a������@3�n5^w��o��PQ���f���ōt�?�s�:HKvf��y�2��M�1�$���ǝq2��qg����W��'lфTӇ���Ss�x��v9�cL>r��/S���W?��Ƕ��C�#�_=�G��;�=(&V�>={#�E¼�=Zb_�L}���UB��j��x��$����6A~�Q��K��ݩg[�dU�Si�9���w,4s�"�������D&�k�μ!�-�'����\ӾE%�.� FG*&�r?o6?��Jv��ު�3A����x��k��{4P?�ߝlm�T��.bF"��:F�L2�:�st�Q]���T)w���@S�T��u*H���//߁^�Ψ�@�b<�e1�>���F5�U��=C����p����+A5���bk���*��⯳�pn��H]۵���N"�;7��dq+Rܫ�6gM*���M�9�s�,�$�A�+�fW�_�-<�?���P��t�C�N�=�a��|�6i���׽�u�m�0>"["͔������Wvg�P=ƽC�L%�%7��G��Z�=��v��v�h�;;)�٤��0�T��C֬������᱁ý]ب�y���_�ɱ�ԯ͒�{�����[+=	���p�%�)����Q{��b{���F����c��&n6w��� AXZ9�]�ܝ^�p�}C}���.���}�$/BE��͊d�� �5ȟ7.ܩ��� Hʼ,��[��[C�-�(�P����QQ�)�G�#�UpqJų��s�����k9mI�^_�]�b�l�iz%h��]���)�BYH�[�X�ZɄ�o�Ou���/�"�"�����3��,��}'�����{`�u5��H}��"�ӽ���%��||��	.�C��	�3?��h`B>� "�5O�;4�����A�iiE��)D1|@�i�=�p�^_������̓[L-4��5�@��F�)���ZKm|3Pf�"�ƟR�q��8��!�V�*�� 9#���G}XQМ>��$j�^K��B�xh}b�g��B=���A�.�����Hi��������_�`���Fk�,��@�#w��c�m��ڴ�7}�2l�׽l�!eفY��$Z�>a��S�w B�nY!禱IY�qNw���c��HM�r��#S{�M��ų�Xj5�t�������Ƹ*��$"���B ��C�#-D��s��߉��h��0h� ��>�R�����>�Ǧ/ u�o+�%C��.�dD6�����ѕ��G��H�(�ٿ*��v�b����l�+R���W7�e�\���OC�>"���([j�|תM��+BN�յy�#�2�Nc���+S��q��0�3oS>�Wz�Ω��'�A�A�K�k��G�����6dۢ�_ H��n�W0�U��<�Ed���@�[��WJ![P����ق-=�����X���U�qd�X�Cg�؞a�}oӾ�;��ˀ7.��
v�t�v|_.�@�=b̆v_LJD:U�����mg��&�O�(��2S��UEEA��n�|���ǳ?I-ͯ/����ۘ}��ez״�ќ�����N4}�J&VH��f���jB���i%�a���4\5�����Y"[E*�V��v�Tr���36��/�����DB������P0�a?Ud	;U�%^��U���d���m�� ~��?i�&d��k��IHĩf���31t�P΀����[�Mb���ČeS�3�ڵ�~�}�4�xa��GbS���Դ��~��b\����QAվ;��Q�5Cu���9o��ۇ���C�~�5G'[����m�H�A���6�瘫!���ؿ�Z&ܸ��?-�B�ߧ���g��>9@���BJ}/3����D/�2�e����U3�f��Z��1^au�gO�i�B.:���[~
��;#�9i�Q!YN��ъ�U(�����K�r�/T�^���)��<���������V��[�����P�$^R�Z�{I@��p��jc1D�t�r�!i�8v�*�y������ït.u�;���!�� ��N�P�"vIqo=_f���qE�wZNI{�$�FP�C��[���y�l�K{=mտ�I���9J�"���G?z��}���Ї
v��2�F��\F�Л�9Ax�l �� ��Dñgg<�KwK���wv_@����n� �HL�c�]3���"���뭂�)}�bEHDo)��[�Ib$����X�uGsbg����<!rd����q�)u0��]w3�8��(�@����#�(w;��9v���Bz����X2;�8��7�6�� ��r n��T7-�˷�
��"U��Gdn,�x�ch"f��{3�>�Y��*}P�3�%���)Q'��JG�*ʢ`�/������M)�K; S,ӿ �a�[�����qo�>��x�A��K�gV��z��G
ެe9�_L>,���E�#����n��o���I�]h���ta}����Y�i�_5� %�ώI��Oj>�8G�=��6����_��C�By-D�6DoY�P��u�`��QԀ�'r��mE)��1����jn;����9|��@�b����3����M�,|�K1N�Gm~s�R�'2^�{�&�Ɋ>���&Z�0�k��t������C�g���G���QŗE�*v*!���ߟP8a�];H�<����섾^;�:$W+K�CzQ�!ȱGn�ʗ݄�vi�����}@�Ї)bh*1�h�����]#��p��1r`O"F�0K�b��ΠfHi2G|�Y�A�D��	Pg��p�����>�]-�Y�~��A����HI�t�9������}�Wq[gS	p�"/J,�k;�u/a��<.���������`1���� ՆNh����<�ne�\���D��C��
J����ں�N�/�v��AoL��LA�|]�R��ϋ�,�JK�j?�N���R�N�:���}W�h�- ye�������< ��m�$'+UYJj�e�=���ߨg��2�A7��R�����G��U ,b4:��A�+A�n� ]���W@S~Hi^�2�
�"��N�hS��2���"NAh4>�u�aS}˺�s:Z�XDN�7�$sq�w��
�Č0ƪ��;EB��"�oD[���leB�c̑�[�:�"�[��������ي8[F��ɐ�����٣mx�d���L����J�_�g�����1Ǆ������LG_-!:#}m"�+i�C��RMx�o5���=�'E�C(�.|�1�yDD6��Z0�����h!k��Mo�"��Q��Fj߷�������9�+�D��}�����e�^2dH�/�q�XW�U�횐�Q��:A�}���ŋBAp��$\���n�X����k�k�1y����"�s�"	�����	%���1�[y��@⛪�v�`�:�s*� �:J�\��s(�IF٪Э�1�#���Dg�1��x�KǄ�g��ԙ��	�I�b�	�-��2<�d�qu���J��ߧ;B�4\����،�!;���g7g�xa���%�_@[��w`^���
��Whji<�U�&#�m�5�&���Y���˼�tH�����!��w�(�뭢
.n����D(@�c�M~����z�c�>�$q��h�� ��	��a�gw�f/hy����$�B]��V����P$�����-_��)���b~��BYȬ�Q&��b�Ɲfs��R)�l�gg�^�����@����~S��=n�I�t[H���ǴP�R���-6K�#ᒋ-��S�i��v|4,~k;���M��6�Y����ce�rip�kT�����2�I���?�~���p2�}��^�Q���N�1-��s�Y늆��e@��{>��|���hN�"�E�bapH��NaL���:V�C�_x�U�^�$�'��!nw$�ЇQ7�J�a͞OJ��4���7���Dy�I�Slc�c�z�	��"�)�DԀl�]��'�����b?֤��O�*Iv�8	:}��\�&[&X�f<0�N���Y\��+��술VWip.�d�9�$��� 2��m9I_��ֲ8T"U��H�Yv��}���n��ͺ�č���$�������
��5b�_���aq)x�W�	���[�;�W[۶�a����(������t��-�
��:#��㡍�$���o�*�{��%�;'���i�V4��>&�h��������	-��e&�Xd�7?[R�V&1��!Z ��Ic5ez�f�u��	�R���j2�]lK#Я	=!\��Q���e~�����T�-\��!U�nף�}�y�qX)T�l��.X�V�4�@YI��4Ў�R+�nuqг�*�@��<V�1�a�KJP`Q�
�cyj>�k=�����~dC����.�A ٴ'���Ss5� �+C�˧r[����9�=�3힕�٘D ��κ�1���j6��ٚc�a�0��2(	1!K�g+ ��èYc�����q�"F6NBʎ�#�h�B�,!�[%/|+/)n[��ɿdAF����j���Xw��]�԰�Q��"|)*����L_��[t��p)�?o6kH��W	���1���ٖ���MS����|���B�QQ9�,R�|��j�g''����_C�m8��˿�Ėm�(튓��m����+�Ti��> ~7q�`0c��]1v��_fz�o���x��9CeT���W&�*���wc�ب�n�e�$f��2]�5���)]K�8�OX�7�r��xh@5q��&j1l����PR<�=O���_k q��B�����Ҋ/���J��q�=coC���kX�4h���0���U�CyK/�5I".vfr�p�X��V6��]��ʷt��|_h�/h[�%�	��آѢ�'�
�	����9���TP!}cU�r?g�B�RY �9�WR����!��i��������'�o��ٿ:��g�0,�,0����~���|N	�yC9{�*�ԝ��w��ƙ����l?yX\��y��H�vA�����`G��o$���a��)g�������^�pZX���+z�q�g�� ����۱ק+���u7����]ö�{�B�X>2bܑ�q>$?]e�<�<g������I�����ߊT��2�+�oj�(�}�����z\R����������K��q�=�A�I�~��*���s���ǪE��}2}����H��#��٧���/�W�r�)��6̵���}V�q�����% �����CJ{��RV��(X����b@#ʏ����F9�:�t����s��W�Ӏ����Y��HG��o��`E �Zz
��pɁqL؁H�ed���D>��򼅡�D�<Gkc��"��*~Η�k^�GI��J�VȂ��H���,����xO�}��������c m�%:6`7����Q6��BA����߃5v�C�~	8��7}i�F+��o�zI�vB�ڜo�XQ�=�;u:m���ӗ�'[�F	X�^�GL1�E���}�>>k~����M�W�2ϵ�tE���đ�Hz�i�:��ev@0HK��qiY��MP��Tx�c�I�ŀ���oǊ��n|_�ϩ�e"�".;�\(S-<m�!�$���h�DG�J�*����nY��K�N���3}͡0��=��D����)�Z��2�%eq�`��>�]0�Q��"���Sp�*��ZŘ��,F�'�ڙ�^i��b^����!,, X���] ��Y�S�;r��n���̵��B&��@jW�.���1�Y�i{��1ot#�~N�>gA��,Y|�k��ޣ�A�F�f�:i�Е���:�:�q߳ϣ�K�5�3�[:D��t��������������vC
擔L�%Z����-���N'�_�♟�Z\�S�� ?�P���	hb�i��������sdd������;���L�j(���gDT�d�%�q	-�����Ľ �1�vΥBS��T�/}{Hy]c�n��=��v#���%����6[>58#�  ڵ~B"�n��g��� �܄c�r,����
C/�pR:�L�V�j��p��V �=V�Ozɺ��C/?��Q��By�\��|ؑ��_R�rYk���b���GS�u����J�_�����_Ĥ�K=�����:ǃƶ��{[��-������Vgق���d��w �$m'�(�����P��d&�*�+ŵ.t���^I�ZUü��5�!�*�A>�U���>�ƅ��U�vLCh�G��)�הּ����9_�۝�8�_�@��u�ݚ���s�}�&�0�k�w��#E�4���_�� ����.w�K*���?��޽=S�aϽ�#�(�թe���Uآ������|~u��ؓ��F(��+0�����a�F�o��cJ^�ǳ�N te�;�g9(��� ��R�b�N.��u?�7�N���C��T���F�k|�r�X1���_�?��"�L�P��*/|,[d%������#p�s��k��D�s�rSÔ�(����7a�Q���לk��%$N,�Ś�r�Gw��!/�Y�i�>��Oճal-��h��\ާnG���#��qk���2s%��;kg��y~�R��&d�+��n�������;~D�6�\0���Gɧ`���ʴ,�����2�A�����9Z�,>��{��w� ���Uh�mK6�P�v�[�Bg�cS<���K{�j,�4/�}��0������cbJ�6q˓"����^/�i;�m�%B�[\� C�XD�a\�݉d�NUܱ2��4یM�ݵ�L���P0��jD�F���Bht���s�0'��v�bwp�qẵ��o�*��Fd���|c�H�u�uF�rvzW�5�YSp#�Z�qXM��?	0V�>Hx��;]Q���A�(��R�~�5^��I�6J"���Ä ���> u'x�Re�[I�C���Z��P��՘�*Ҕ��2�u-y�7ETR��D�����b!
�}�a:�9���@
�D���m���=yM�^�0>�lϽul���^�B�ږ��iC]��wE�Uz��Q��5�S�g�������n^���)��"b�N��cY͊�
0��k��/o�̉�9Y�L3��L�W�|}��I9�-Ő�������M>�n� �
L�y�O�d����e�Pt��S`����>��F�	��*'v`%�k���#<Y(e T��:!.]��{�v���굜��|�\{��	m.��$�1Y�e3r
򢏶�N�Z�t����0²���%G#f�v��_�*�$.ޞ�s����ZMŔ���f�l�?6�{?��p�U0����B3�#TUD��l�>����� ���s (�8.��%
YZ���4z̟�=��-it��`���ANA���J������Z�!�^G�|E>�J{�q%�F=�sX��a�3���ǯ DWT��}h2����8C�f�X�g���A`��=l��8�ȫH�����L������Z������@��ǆ)�,K�E�zU��
���r�f�WP���Mڅ�*�9����t5��#�t���X�� ;7�oӶ�j��B����#��7�ƃ�X݂���(B~CVR�����=����JnFO��?/y� �=�W����I��)hu�4�[�K�m��r�{Z�HM�$����$���e��.s�\˰��Z_@Y7@�����-�(�,�Ro���ۼ��T+��G�{d���]�xzv����8Q�A��}cX>�H��OO�Ee�6E"�67���	Nw�~�ٵYKG޶���iA�ǬU���e��\�b�?�X!5�VFl�S��_p;8�O=IK���l2\-#V��Tƥ�:�rtb�^q \�l��s�0C^�Z��J{� ?�"�$=���7��77Zo�U�I��+ϮC�M��a�k�6J�������-�,u>�"pE�	�H�۠¥h�,���v�qG��`�iU�~î�"��s�ۦ�8ϕB�5X�Z'����jϞ����J@S���"��S�������@ˌ������[ȋLg�:M��u��a��d�Kk���6`]��3����	X�Ut�_���]X�����7�4��#:��n98L(j�Ű���M��5�����Z�w�A��bh��5�!	o��yެ(m�� �1�S�8�$�1UB�(� G@�ܫ�ո0��;��,�h�dT+>J�L!���C6�ѭ>K�*r��`���b%�<I�\�/�����s�'NQ� �3z�38��=ӣ���oM�%?l��+��Kڏ=,ԗ�fls0l��g�lw��_ �v��
"�Zy��b���,��r�6q�p�n��� q#�Ǧ�xWeӱ,`����aRt���z�Ei�w�1!e(V P�t�Z;�ah��Ҽo5~FL��l�P
���Z��t�W6�$/㈶3��D���Y��`2��r��|���=J(�f��i�m�B���ew�+p-xN����4y\��+kV1��(��6l�*��+��Z��6;X�H��Kx�<G!n�B��2aW1]�v�1]q[�a�D5G��Ɉ�9��ĥ6�{��)�˺�� �����'<a������>f�i!D�L+��®��ԝt(/�Gsn� �'���7� B�3��e��2���uu�o��Ob�pki���CQ�Od�b�viN�ͺ�;�/+��;�_Z���u�H���܀��]���Q��#�f�j�[�3����8U˸�u�'S�
o�7�� xӻS�}��G��"q}�O���_<�,D��Łg�踞蘾���k�]E����*pbE>PZ &�bF�����<��FN�8M7�`u��hX�N�r���xpp�Yaǯ�=�Il{{o��cS�k�)öp��>��:�)�<�Vo4�s^A�!&n����{��AR.���b��94��/�
�w���յy@��B����^ML� ��kN3N?���0I<�L䖡��pc�+ ��k�W\m��еelE��Z^IP�XWoPRr�������#ׅ?�f���v�'����B�q�Y����7��W'���@;�w��.'G�s�j�E��4T���mi���[�d�1e[���~�j(K`W'�����?�j�@��!T��]d���gk�E��I]F���MJ:��o�`Ϧ+M�WQDg�7H��� +{v�i�8��]z��QE�b��ם�E�~x�[ �q��<�=���L�fY�7���}�t 
A�:A�-h����RM�B8�����}̔�%R���<��"Vܯ$x�1t�@ē^d`6��L�7|~W�V^���Ěݎ?Nu�� W�b�����"��
�g/����W����_?��Z���<��+���xqR-��v�����*aZ<N ��|VM+�w�� �Z;�Xc�%>����d�yu�k�|��/������3ٛ����=�g�GD����KB'l��y������d��^p!v��9��c���y��Y�
�&�=�RaGr�"$=׃S:ғ����>
L_�)�U1�W�m�<n����1'��%����$�������c�M�J�G�L�IOF]S�s�Վ�ή�C_����Z��NH�	� ,Y}�~.�w>
�haς-U�_ۣ�E׼a��3��P��D]dz������	<��W-�}O���ٺ�ū�����v;���.��M�j�G��z��p���vKH�����̈́6!H��rt��g����>e��!�{n=�jj	����Y�z�ќ_�Ni���l��I�w>6���f�޶�a	Y��{@��ݖ���oK���w������h�<~-ZZ'~��Ǐ#�1�r\˥7E%�]�r0�۹M���Y����r� N�z_Z���՘�*�+��!��M�u�.�fԿ��G�U\d�p�P�r'��������O���9�Z{�p8�u7��x���0���5�ϰ�B�ݿ���wuH)�6�a������٢G�mԨ.�kB���J,e`	�5�,�;z#0^�G%�YX��)��]�����vAX�Y��e�0��F�V22c�Pq�:Kg��+2�����#���G�O��'���?F�8�G*)Pn����%�qv>�-�lz�ױ�u��9v�h���tٍ��C߉�r�[�������v�\��35HB;
����>�ȹ {�kŁ�7d�>d��T	��T��$]ϓ۩�;/��p��WæWS�zm�"�$S>Q%B���_Ѵ�9��C"%Z� w`�ԡ�o�ߗ�&E�岅��	��2��JZ���*_�����;^���"�.�Vr�ʛ��"���>�	��8������P�@o���O�#:��!�7,t�ΣL�Đ*(�Q&*�����j�1?�/����t��<�`����`�!9]���E���y�G��oDy��xJ>�v{%�c���`3RZ�����c#{Q+��]�~��%ܒ�v��ݏ��n�T�B�^���p3�
K��2�v��V��d�)&���ծpA==�G?�
�sC��i��T��F>Z��NΆاr�=W[3���m��:a9vň�E�i�0�Mc��u[����ʽP�*�XM:�Pk�-���_�8E"w\��B�F*�n���b�!w�l�=�����w*b�ekD�B��|[��ey�E|M)8��7�G*�BDʨ��ĭ<���?�
F���p�*��k+�)St�U��t:|(�6��m)�O��E��Q+��o�H���\�����a]vkv.���W��n�危S��>�B�����F�%5�*��j�v�˳G�(��$E��P��0+{�Z��H�~5dϖ,��V@Tv?�v9}��UK�~�X�F�H�0��V���2Yb��*�#��@�:�_�Rx��^��7t������j��0|[��:���BC�evxʦ�D�r��� 6���kR��k"�ބ�M�������E�ŧk2��8Ŭ���6���\N.e6�D���[������u�\|E+�>��*o�V�k#s�8��WQ;�i�}h���j��\����s�UX*MT�ԿVm�rσ��1h���|�R�lz�G�F0��R]��ȴ��U#� sM�l����ل�2�~Z1�w0��T_��2g���8���(Ε;* *��_�.�jhR���D	��Ƌ��SX4����!�݈�=�c��#���y��S��k�}[�`O�>����!�=��W`N?��h��H/��V�Q�����Z"�ҥA �%/�|����A�x=�Y���^Z�zB��ZQE���d�#n��L~S����*T1t�ȼ��^��,��r,>?3q�ݧ4@����1���C�Ae��q�^����z>���~֛@�A�t��?�
DM�_ԙ�G�\�P��u�dg��m���óS��"��+d@��j?5�������˝������I��=�5a��2n��E��L�I��]u�W1�&m�ބQ���ա��R�Ϩ0���{�Ǭ$>(!��Я�Ɂt�O�<���.ZN�ui�5�::4LƆ���M/6i�`��s�u>��,ۯ����M:�N��W�`v!�К�8���Kat�ϣ� ,Z�~Ls�P��Dj��T�$��U��*}�As.���dI��hP�0�nx̝�V��$�bi��i�'�,�H@\�2��BhC��9�QjW[nqA�g������Ꝇ����m���Ra���y�":Ʉ�����3�a�y�ʽ�X/Q�n��b�sxD�P#�H4p�_���?��Ը�W���9����˭�)�T{�Q��N�4.x|�� �����Z�m14�炦�3 �J]�����(CŰ�=��]�V��;
�'΍���L��aE��(�ě��5?������j]fTk]�׸�M���N�����霿�X~�H�]�b��P�Y���$SP|�r4�2�[V�Q��[��܃|�7���P-������3��V�%�I�[0r�"-py�0�Gh�?Sm�(Ug ��1����þ���P�8S|I"��N��tS��:�j��{ R�~+K��]�n�ވ������7��Y���8O��"ﱘ��#u�<��Dܳ[�.���mmQ�;���\r�@B!��8�rV��[�|��|"�����5e؂s�S�m��	��܅j'�u��� 0�mo2.�l?���Q0��ћ/��rў��|�f�ݘgg)����~r�'h���kv�/��>����Rn^w'lL�:�G�ێ�g
��0)p�ͣǒ��ۼ:a!ʵw��M�<���$`��̻���ǜ�DfQ��Z@b4���焪�]y/���6�~᷅��0����Y����.�������aM�q�0���� AB���Fi%�%���"�5L@EEZ@@@B�ѣk�tw�Rb�6z4�k����7�q�Rw���'��y�, �A�'�d� 0��Euef3�ۏT��5x+�2_S�7�X�}77Wv�+���ϣ��8� ;TZ�r[�!�D�ʠ= �Q�����߂p'�޲BZ.�bCG�30ۖӖ9�ؚEb�j��F��	Z'ʅEG�8V{r7�O�W��We�Ǎ�O屚����p'Un�7Xi�u���Q(���
�n��&�}����b���h�?Ka�N��a��ɲ�5U~'Z��׻����M%��`L����見�pt#����ʏ����;�:�׈�Z��'��fO���1֨d������,�/��E��䷟cq���9�8�N���,��,�����7l���:�.P�f�S��ɗ��Hl=����G\	�x��a[�����?*#E]G��.�l���4�� �C��W����Z��y��G��.��.I�olZ�H����p�N#�c4QX���7(������P��667Q);4�I2�h���f(Z��5N����OI�f[y�����/m/]Z�"d7��4��$�7�E�<W�!o����G&�Y��]Eڣ�H���7�����2��+�V|�|N{(c]I'[GL��)���4l7��F}Ĳ|s���ϟɸ���7|�o��m�njT�ʋ��<$�xs�� K�2�{YIe�Η��r\PJ��G�t0�0i���\��%kv�9����b%��c b9�،ryA'{����͚-��[�N����R��]'�@f�vK��b��Ǥ�2о����ą	^�e	+����nE�v��$�6���V�����E����ƼT�У.��4�u���:[1�������C�㐛[^|�!H�)'G�E$�D.�����Yo������'�hRq(�.����鱣�q���\[6 H5/��Z{���6���@���PP�ˮ�~��Nt^̈���/���=�n��Y��L����ו�*yͥ�;�p�y��6��}��45�²�O�����]w�}����x6�Fk�����0+�L��i���h�}L?��4�i���V]ǀ|I���� Y����&&���noQ�)��x.]��ktj\K�:�g3�%�v( �~[��#y��	!�z/i�u-(7;��d8��8������;�׮_�c@9t��k��au~  ��_�~�&�/���F+�C�c _3��JqG��x���߻ͼ2���H/|y�	qy��zM�ʬ�	Er
k�e��N�'�iZu��S҄R�ٵI;\m����\�-����}(@%dc�R%��u�B����2Gj���/��O��R�2=����7�Q<�l��d>��n��I��[�� O�u�P]_bh34�N�s�'����w�Ls��a�Z�M.+�*�qV
1a��:�܉4��
@��jpWN����e������{Y.�I������ķ��@ꉓ���\j�N�ЩsKg�$[b�L*��P�����Q*�
ͩ�+�G�,�V�[WkU�F����z �Y�I��1E_$���X�9^�S��gRW� �%�H%dw�NG�,���O
��/g�2���y���h�P8�(��7�me���<����P�/ܽ�_�o54ЧW3n��������)R�߈!�CFA���X7N�5~
>2���/]A�N�Gw�m\����}ƙ�Hż���M9�mE��<Ù���%�n���]�z
�y�?d��u)N����p&�H/������a���;�o@��m�^0=���\`G
 �|hN�o� \3YQ,6��8�s�c$脸���@ƥ01I��^�0hԜ�X( í{�y�t�g��d_q��e����M�:�- �K�`�s��-N �d���Yp���]�����j��%>z�۔�@�_�&y��}��o��k֌���(���L&Q:���b��0�A���r���
��o�o��`s+�B�2�ʬH4���}�Υ����z!�e�����[�[��"���1����o蚵[I�N�R۝�n��e�R�Ӷ�X�tY1�ת�nf.҅%��v?����$^��L �� &@�̐�����*o��<�cJ�$�C��<�sA��`ho��)�ad��(B����-Z�13�> dv�_<Ox�OpA�
��3��]�a-�&��1%nya���\v���m��r�kYe�M��0�y\�ύ��=> ^��	hMO���z|��&�oIsV���>� 4$�FJR4��x̴8an�×�s6��AfO��Aqg������9:��z�T�$P�u��t9Ώ��i���Օ������a<]��ZW���K�L_s>����n,i��M��ҁ�[g_EB�_~&0�ˬqZצּjM�W����Fꦻo��~�:��ښ̳GF�C-{��A��?����X��xI
����2�K��ޱ/#�8+��B3�NB�4d�{��HU�C����z��	!��v�E@�(_{7q}��}nӷV��^��7�|�Lז-��4AML��3b��f�1V���s��Լ��d���,+�S1�I�p^_����+�c6X����GI���W ��c�71Z��q�|�0h�G�lÛBY����4^.e]����z��,�='��5Kb֢E���+~�Q�b�)�|Ҕ! 
�*6#��<=��X��i��9H��d��T�Q�����9����*��N�e��U`~��L�+������*t�x5l����]R�l��@Z�+�M����#%GW x��Բ������� ֽ$��"]���]0nkd����qYDcn�Ƃ��q��\ ����)�YUs���	��ly��^w�3Δ4�j�T�&�s'�L�f<5����,Ǿl���i�Ahn�[�ڭ)����.L�H[��5�/tfveo��Z��rqq�C���/2����3�:lv��!ɘ?��:C�
�t��d#76��'TCUR�N��Q��ܺ���餙R�6�֔17��ַ���P�%�M���inO���{�ي���'���	��3#����1V������0����2	��������O��˼(|�犙]F�m�ǖ�+���9�B��/�e��Y�.夏Q�vɯ����<�VwҒs�!�z� �]�ԯo�x�h-�[^a-q�4˚�on�ѧ����P�t�5��Z��&��g�Vb�G�FO̙��nY�v�Z�.�_�������q[]�%ճ���O-:� 43M�b�'����/4�%	��cc:��WF�i*H�п
�Rn�����?UX�I��S$%&��ݚ������<��;Ah�"� ْ��9�ka��ܠvw�)3{p�~�B�1�t���lI(`<���_m�Xr&2$:��-�A�zG�k֓0�<�Қ7G8N�%��lW`�ޙX(��H@�6�kP�j8��wRdtZ�ʺ�i��������%!R��idM��g�r{fۊ%1P�[�����V��c�VZݭ�e�����r0Г��y�hٽ����?t9<>��������GV��A8&0�[����`�j����볇<"�p{I�J ���g3�u&��������G�L��	��JV瀄�$zT�5��ޤ�E;�����K@�ON��`���AzP��q�c���}�W|���_|Z�1 �]���S�LFV�vT.J��o+����V�c�������-J}� ��2���-$?&�I� ܬ\���>�B�}�I�N���۽po�y�h��-��V��Qn��꜅R�#�+�ݠ���En��#b��K�����Zw�f��}cWrK�/D7k�(���[ķ���c���#��$��8:�N�X�LB��b�D`r�=�_�4=���̍�����w�\��].�100�E�i��J󅹢^Ӣ�c����=�,��m%��Vp(��xR��֒���OzY̋b�O�K+��|����t'4���*n� ��=n!���0�����(.Sq�S/���ˇ|�PXZ�d�k&��[�oہ-�5�~%��sY��� ��đ1�Wn9�F/t�j��F�����R�i���s-���0,��2�V��6�-Fiq��_����m5sE\g�D�eךq[�r��`MG��X�}#P����*��ԅ�Sr���*W�i��Cӳ� z�_`�}�PC�I�h��`.tz+�|��|��3?�F\/�(���}��������
jfQ	(%e�*�m��?(��@�$��Om�g�7j��u
��Gz.=�ta|2.P��v�Ί��::����"� �01�]g���R<����f�i�}+� ��W�	?3ӜXny�	�n�v�<��R$�"[<���x�W߲)�7����ʼN��7'L��H�]OY��;�Q�$hm�~�o��R�n/ǩb���]KD����%�~���ߐ��^��~��j%��Y���ڙ�ė^�Jѩ��A��Z�L#�$��w�C�;�$��8���x�h�-C�	Cͻ�����4> ����ٿ�����Y��म��e�󻓔I��i�8z�~��f_tLzϗb a�v��+���]��1+�s��6V���V@Q�-��<�ԣl]�|P��������B&[��%M+X:;;��O�<��E�z�,Eʿ�O<,��w�\(Π�[=�� �[�m�?����Y���k����n�G�}( aK�?���,2�Md�/
�o��&6,��X����(l�L�SYэ��h#�S��&}%B.漐�ч� ��O�[��ԯ2Q���OS��,���J�A�&�'+p�BbR(�>� ����|��$�\�m��x
�Q�,;ܷ�������j��c0d�l &�eg����l�s�^�l�d!��(�����5��U;2�H�FT��F�!O���-�WʝA#G�d��H�����B�WY����4�.��`=�d�="�y�*����$~<�Vd:ώLV�!��xb,��Mn������1'L��Q=L�9�דϱڑ�n*ja�a&=�_+4�.P$L��1%�	���5 
+��Y�l?2&�J]����ղ�;H��2wR�l�����X���� �������U� ��]�K�b��j�R� �O�fP�BHsJ��
˫p}*��C?d%���ߚ41��v
��w��	��B0� ����[5�V�)T-��
�w��K�eOG��$7�JT�ʚ�
J�YQ��ٹ�>���ϧ��]��q���}]�0�S�&ѽW���Ʀ�ye��DJ*7�a��߹݉�	��G����(�0�դ˖+/�@s*:���o)�X�'���bo�=�e]z֜�h�]����ų�R�Ν [y�F�pO�í;������;*6&r)X]6\�~��"&��ɭ[�f���ZsK1@��\$�٣%��t.��S��-�P5��*D������|�q5��z���<Lq���ۿ1Z2����?{��??��?��?m�3���?��&�O���w09go���vU����Z�4@1��^8���C�kd�M�hosJzdԴ�h��פ�v��"���8u#~I�'���7ˣ���Q�وl8w\�Q�	Wb�kk�q*�*�IqR�Å�O�8�i��w
��"�z ���t�E���zᵄ�BiW�|T�l\*S�����^|zv`�)�I:D��lF�Ccc��FY�D	���N���7~�a�¼��P�|
#`H��y/I���g�&��/�1O؇%��{��&󌢓dqO��wjaX�2.+���q�u c>��}��MGHOO���B^���	�F]�6��?P~���ˏ�}������������ū�/���*̈j��N�;��S5��Wi�U�h�I����%��)o$�X�'����x�^�Nj����6�Nw�;���wڼ�o�!�e�R	R�/�	zY�P��3<�Mi��5?v����J@o�\����&���n���K]��yi�w�s��Gȩ�����xj�n:	����Q�������!�ĽB���e�WuL��C����ֈ�M���Z�ư�H4�@�b�hg���g8ū��~7�V��^-#������Y#��J����q�$�:5�'z��nyL�yV�s���.�����<!�MW�I�q�g}%^�l_�65?!m)&t��=�5�^�ЉH���|9z8}��!Y��i||����㥕�+>����
�|��Ǭ��Fg���$ŉ��M��d�Kj��(���d�	�_��߇�+��xi]�5��������'h����mi/����;+E:����;d6}�s�XB���X���ǅm'�2�ʘ��5"��>�2��5�]S]k��V
�ʖ����G��<n�?{�z}6H��m����^!�v:�r^z��6kz��o{f����������Z��uf}�{�n�eXn&wSg�ɬ�-�����ߛ�U�m�Bb� �q��VW���0���)���_B����Q�l��_W6��B���^�\�@ؘ)�-���TM����]5a��g���¢�?�������4F�g4����;�3�s�2�F��0�M29���p��g���d#	L0
�ZJ�z�v�(�m-�](I�(]d��I?�y�ڨ�s+������r}J/��`
_�Fڳ���Ò�C��9'OFݪ:_O.�u�w����k��Ĉ�wk�B�n��j]�`܍�移����(������JF�\i���1Lպ/j'�G�H� �R�jXu�G�pPP��x�&U3Y�/��~�Y3	�Ǩ�.��5@���}n�RQR=�X5"���M���afzz�*G�^<�me��w�dWݎސ�C|�;�����F'Ů{�0��w�O����?l+��ZcËC�mO��Ƕi>���A�mY!��^c%Y���C����;�S��پen�\	��H�閑�;Y_J2�X���E��TG��#\������V[D���a-�&�m5g���u�O����
ɓ�x�y��N��Y�Ě%��n�|��ɕ(��� ?���*&Щ�>c��N}���~%>~�A�vy�i�	�L5�������'����YbM���\��XEe0�@�銕�I�Y���"�$<ݵ"F0 ��_����R�
�tEFDn>��f�M�L=M=�_�'į�@u���"���vv;+�&�`��Q���/�h�>!�7���Ք��ƣ*�����s�Qq<��%�U���1];2?����s=3ٻr�qn�(;���n��DH���m��"�:L=�0������w61"�-�����Jt����������8��d;<����~��i�Kn9Ϟ�[[~�ͻ��@Y�:it���D����'�:N6kw���
� P-
����w���io<�� DD��s�J�n���,��R�A?">n�����w.��9��?�S�/H��Y;Eo��ڌ���H �	���'��%��*++M���`=��`o���u��TF㶐0���Vꑗ���9)U�C�^ 㝰�ۢ35�W����9Hk�d�AO�B/��s�n=m�/j��mc��/�M�2u�\]���N��R=�Y�h?}��&v<�����x�N�.���hJ5f�/o�Z=� ���BM����z!J51i;!ȎeQ+���zi�CާGĒ�(F2���4D`�t˱!���З���|�3SU4B�t���w��K� d�nVڣ/�.{i��5	��K:���H�u4�x�n􎽛����O<��Y����=|�Ϧ|+���
��O��b�gC���-�9@��U7I�R�Y(� �^����!��䯺P�e�y\S�%�x�G<��8�zlydtnEd�&�4��T53 k�e5'>䓥�>�c����ǈ��e��V������m������^P�M���_f�a��1�ⰶ_�Ny]��L6r���ن<G;?|ć� n�`nЍ�~�頋�I.�+C���l��R�pPf�������g��<5'I2'
�c�)an�Ӝ����pW�b��~YV�<��2O��z&?��S�єQC-�CL�N�W[LXf`
����߈��>��&�N�ƒ�"�*�HD��%4���'-��o"��yOޢ���@��2qj����Ù�Bi�h�Zb6Y�sB�	@�����U���,���dW�R6Ά��P��7T��;�,=�I'�ꏭgl'3��ݺ�����WHYs��[��a��@��Eܼ4��{c�	�+�M��cN'��y�&u�%-�����Y�{ߊ�Y�{k����8^�o�=�A6�CT�d���P�7:s���
!��	���1ʐxu���X���9��wyו��*�6~������꟝�.s��G�\1:0� ��E�	��Ց$�	�0�2�����ɔX���6x�q����	UF��%�8������W�Wq.-W�Y����>�g�P���] w��>,��.�v�RU9�_��{��� �x`P���Bwc���P!_^R���]��k!�nrSD��*�=���.O>��߉�Ъ�6�L���۴BJ�-�%�m� �Z�T�5R���P��݈NU
P�T䇄>�	ںR@H"zq�^�č� \�>����^e�1+c��XK��#}� iXR��G3�V
MO�f��z�T'u��Ub�U��ah����bdp�D�b��@��'��R����C�O�5s���۾��|�c��}��j��6(�q)BT��+�+ �:�^V}S���7��$�G��ɞ�7�n��W�z�7j_��@(�6K{w�|�M��B�u��Tc+�d��v����r�<U�$�Di�׾��
����[��z�\��7i#3k�2|u�7� �@:��[wI�D�N�Ƿ(��ijNq�v�s�vh������W-����}�+׋ee�T���8�=y:�wFgFw�yK#�-�F����ǋO|�~��V�[,Õ!\�U�;/֙�@eWg� �}u���|���T0A]�����I�3��SE�n����b ���@�N/��Rq���A����^��j��8��H�1j���ݕd�fę�!^�H�%������a!,�#4ޏ`=��v���IW���[��|��4M�%�+S�թ	���7���>�H��z�'�7T�z�����-�(}F�N=��1��r�����-O��t<���v��p�LH0&�'��rמ����Z3�)�Qٻ���x��ʟ��q�d�K�>�i�5kO<�ȯ6u���{|�a��R�Nl��n�S+��@�N���� ��� ���Pҝ���ϐsX^yJEJw���.<�V3�:<a-C���U�Yȹ�S��י��vׯF�����<�N���W|�+��^P�J�����8{���r������ZAI-3��#<C��`r�tsep��O�p����)�BvFi�# q�H���i��h8YŠ��@?,ئ����_h4���u18h���d��r�)(e��8lU�9Z�H�}�WOl@=��|��������z!"ǳ�2t���P�T�k�v�B~��Y�ϗ����������(z��g�<�K�Od3��%�E��d��*_˜(���J��&Օ�OL����+���}�Le&��^��M��a� u Y7�����ȉ%U��W� R$�����-8�0���~d1ډ�X���.O�SQM{���}�CeH�ih�\���+����L;���g/�į�D��ao_�f�aK���������;m	<W"L���Vl��eK���[%iA�^��c#�4��B5f�L�r�� ���Xa�
���>��z��6_�r��hT%?�w.(��+�����[,�b~�Qf/�S��2{�l���XP������s�lQ9��ʿ���b���Uk�<>A͐hߕAٺ�3���X�V15OK��v�e�|7l��!���]Q��e��q�#��h/I�(
�ʳ��v8h7�&뾵��M��m��ҩ[O��%>�}c6)\���ڇ�o(�� J��ԇ�[��i��;P0���������fa�t����������z>�H*xĳ�
v�}����t�U1�ʛ(r���ؙg��2��<�4���w��C ��4������ظ?h�v��{6����q�t� �v�>��=o������pB��V�L�(Q��0���-m
�!T����<��K�M�3�s*_����ٽYI��+�h�-��>e"���!�
H�+$>$�G�*��$�2�3mJD�	P*z�D+��~wSs(2Ll\�Ob��o%����T��^�[N����):�#t&rC�k�y8��l�!i�,X���jl�p�:���/⥬W�֕&�]92�WH���С�������ʯ��1��fz��Gt�a���d���td<w'SN�-e��쫓��+c���0�?�́�?u�B���6Iv~�)<�b(.\���7}G��J$x�Q�4���͌+�v|��A����l���<1͸}�T�2��F�ke
 � �"���6��W�r�V�����~,�vZA���T���㇃?��գ%y��+V^>�-����H���Iq��a6���i׈8���rDs.Q f"Av�~�9�b��Y��R���� �D�d�i����^6�ꇜ_�Ĵ(��V�V]!���ʀ\�M�n
�<,��w#aBs��"�Sd�V���۫��<��!j��D���Uuԭ�k�:ϖ�F����]�Qv�/ʎ��Y��е_����'�d���p�ԕ���� -���}��RR1�r��z	���WH�!nᬺV��E$��sd��t2�����	$ͧ�'�����O���y��N���q�YߍY�&r���*�	��;�Hx�����XH�1�h��=��74��D=\����ưNȄ0K�Uu�$%�g��_)�T�fci8�E*�m��:��c,�^�PhLa���l��W9?�?�����2�8.?������ WNX�:E�W#2�Iyf��-`���8�Q���(��"'d;�.��ʍ�	�R'�P-Dq��7���6�ֲg|�t�����:.k�������z����"ɉ��S�u�5���^Z�Ffĩ���^�./��ҷ��M��H.�h|��0v/����F�j�.�����E���G�#����M"��J���B���qj��r�[�谄������'�5F�]�����>d���wo��6��u��z�M�@K��9�s�f����\D̘hqg*x�ü��Nd��P�n&��`�<�
��+Xq:�zY��U�؄GX�ˡߑ�+߈h���,J���f�1'F�Gx�H�Y��r���3������_�qs�t��o���RǠ�����G����Xm7�)���ߡA9M�h	,c���	4~�8���2��y��� `PV#���ZE �E����_�M#Mhq�1݈�����i~��$�,�!�j�����9_� ������y_�h�FG]�~Y�3�0J�=�7�q �'Y���W$������8�q%�0=�fPV�P����&��>��̚�iɛ|�W 'f�%/��V��0�g� �C��u1]P��ЗC���&�|ǹd�	w��Ɍ��xc'ٷ�>�0|z0*;sXu�������GXPX�8�e�i�]>9Rm�>(3!���{(UB�VJVMh��|��Ç
���7�����ml'��F���Ѷ�7�mT�"ؙ��p��O=�"�-�H���&��ec#��������?خ6�^F��6�9��4b&-	��>�$M�<����=rCf�P�FW�������p�c�����K�|	�}C?�"����y��PR�u"����?C�?C0
҉�d����un����{�-	�x�����o������%���9�q�p�9�i��'k��҂�s ]��H��% �چ�嗨��i*:�[��O��z��H}��a&�L%]iIW�*i`���]��Po��W)r�R�����d�a�}iO1��])E�����ϴf:�H�ry�iY�PԼ�gm���T�H-�z}�)�LW�Bv���4E��	@��"�*��_�.�����Y�aL���#��.f��9 �􎶰�T5q���! ���̵�U��Ab��: a�N={8G�Ӳ���*����e#��E���{}P~2x�}d/�4�-�,g;ԨR��]z��H�^�O�[C9s��N�}u��J�}Cƨ��UqiO%j� :f���0ᨤ�I�f��.)��%	e+m�i�Co�R~�涍s�8�S���dj�v�����Θ����W�N������D&�2v�Y�8�;�2{&63
�I�D���2��儐�,>�_G��9�z�k_F>�Q�.jk6T�,?��>c(���L�8
�E�b��ρe��/��;L�6w�15� �l����d��h��Glh/%:���;�k]Pk�eq�\|�'f�֦��iS0�����Ę�F� F�BT{����C����k�����і:��o�~.��\����0(���)<<:�UBڼ���C8�#v|u��h&6ˁ)�S�śo2���6����� Z}�r��mc��__	���G�_dN���cX�+'kj�B�ڹ�qҐ��C�p*�W���wM�*z?gWV� c�mm�Z�5:
8�`9�(�:B^Nc��]�C�Z��/e,S{�S�$f��oq��t'��Y@OǨgY֦�;�N﷟1�-3�+`<?5ew5���f{Y`�u]?}�*D٤7j2{����4�p_ٟ�^�T3������
�����b6뙏Y��LJ��E����?�*�ݰI�.��>|gӹ���3,b���A��"�W��?�l��nuў?�9�i���?i=��8kM黤`%�4�
� ѐ��#
���v���O㏗���L�,��lM�A�����>sIU��@!�*N)�j�6�(��Pl�I��į�u������̚:���A���K|��nj4����׾�����~��?��r�,8����Ė�%ę�R�v�����#�k�]�Z	����ᙡ5ΓP����D�ӧK��ok,|���#@oӎ 'X�Ϛ���t;�T�̗���l��$�#�+=�0�f6H��U�R�e# �������tm���q��X��v8c.�0�Q����Y�)&�*��i�XFY17ђW(�Z��{���Ͽ"f[{Qa����^4����V?�D�Tu���l�S�U��A���=#D~J�,��ĝ*���uL�'v�5{�1v8�'E �й2�<�)"b�m��ܲ;A�M6��Ӄ���u�d��b8��$A���P�u�$Rg�/z��Qy��sx���� t3�X4W��@ar.@넕-�G��o����N�+$��W��Ye;\O��`ɨ8���{�6V
�{���8��V�� E��8��4p��䥯*���CV�x���ȏ@�}pn�|�9��u?I�&]�BElCc΋Qb�Ү�u�{ŭDa�7�`@��������λ
 )���,��_
*7�����5�b-���ں�qGEO"#��h ���Zό��{��딕��.��5���kVg4x_!��$E�v.]v��
�+y��
����g����k$�e���Ws5���k���K��4x�P�ə�<�H��Gbq*zZ�9<ľՋqTW�ШBN}12Z�G|��k {�wՇK� �KC�m(V�/�7�n��ns�q.���d���x�=-��hd]�����d��h�B�zl����ߴ����8�Ei������ͭ,GR�)e�xU�N�mnOx�FoۮM�02�ڋWr�'�4��Īg��ǟ%rnZ��`�I�C��E7�9a͇���2����b/��ل+�~�Ò���"�}1���HB��U'�تP*56���d(��r��&�q'8/#u�\���g�$�D=�AD4�&57�3���s���w5o}S�90����P��*%�m�k||��&��L��|G����x묦���}��tz-ũ��oT�@�1�<0=�2u�S>�,�	4-���辚��%��,G�Q�(���t}�*&��P뗑�I���ȅ���u$���p< g��[&8�,� �O��7#�{u��)yr���\��C0>����{om����*��
���+�%߉��'�8���-+�]= z7R����ɑ?z�}h��n�k�^�u+gHeϳ�J��jL�ρR�&w����}9>���)��9'ǽ�Υ�R��>S���,/��q嶭l����ݭ���f�����
{8��?#����{�d_pŨm��S>V] ������"�J��cb���d��O���ΚAIra�a�E���犉^�.HS���7�+���*�p�;��ʦ�g�Z�j���',�T�K|ީ�|A�2�I�y��OVYV�o"y��X[�IQ���c0%��U2�����N%7M$�����j�9$��Ӳ���J�1I��\� JC*~'p&�"\:2�L=}�l����o�Wxޕc7��+�}j	�����g�W�9z�)�M�c?��.�� 7����.Cw����LO�|�����ܹ�*78�;(��=��;0�I���d�@��d�X���Aꮌ.�.j2�%ŖQOCC�Քr����� ����0�׺,����F�t��'�:�Qa�li��|H=[�v�T�9^F�Y����jH`sV�zye�c���*L�{K���zh�a��y�b�xpHg����ͨ[�{F�,��խ��S��P�X����j.�b :ޕ�φYj�� u[#\���]5�ȑ���n���<�绘��g3z��ң��
i�
�H����^��w.ֻ.��/��G����p �U����$�ϡ�W��`�+SoDdݴ�q�����᫰b�����{�,\���_�>ջ�\�4Wյ���[@Iߡ�2](y��+�kiڴ�:�Z/�?��gW��;��T�6���I�Cl^������X�x����E 7#*Y&�OZ��U[��$��·gd,m��C3�8��:n��hEѠzfh/,+>>Y��c��Gyk���z��q\`5���7]Wt�=L�]��%��@N�!����=� �J����^�Q����صci�����X�xE��m���2��TRt����hK~�S~��UMܯ�]����螺����NWO~8��u�{��o��BX�zf���%�J���6�����_�p�W��#w5.h�}���������j�XtWᄍv���n�ᱵ}��E_��?15��>4��������V�M8JKS������m��O�]TN��C�'��s>��M"�b��������ꌖ�e=7����-��5+4�1��}<f��`��n$�B��l�^�X�PYR�g
�6U���Do��5���W��ڼ�w&�U>� A��~J�g��H���%ʳ(+�l3�ҝ��y.�P���F���2S�sk�����W���J]㓜jL�*���+oM���O&]F?�|ĕ:8d�g�hQV����FU��m�tE{�gB�?ݾ�Jį�Uf���i
��;N�v��̥���YN�x����s�ak��[['��}_��z+z����wu��SD|.��<]p���/��It_,@��̕��l��`&Α��a"O���m�}arj�@7a�����)!Q�]��M�M(*�����k CtE�z'�(v|�]�-�(%b{�U�T�aCA#/���7��+����%�lĸ�ɍ�v��_������.
���^~�f��7��_�����J�(�/�ư����Bw�����2 K��_���bF�F^x���\�({~ȩ��7
��)�66�o���W	7��NU��
��^Z�Fr���e��]Y�^Y����:��F	HWW��Z$Tu�kVV��dn�xG�r�LL�=���K�f9&��䝏p?2;\�d���d�Z,���EiJ�$��+�E���-z�鳍�	=��+����f��;�W���W��j��=��Pe�"�ᔯ�F~R48e$�����*_QO���4j �iG�UΨy�7e�� ��]��d�*F
�C��\.ZY����3���[53W廬�0��8�Α��쵤w�"= �'�Q�n@�h�p���Y,W����G��z�L!ȫ���t.�Ͽ���!�k. :E��U�7_ T�����P��6�ࡤ�b�W~CI���K�������t��X�K<��\54U ��ި�{:;�T��X�,g�d"{!��O���^R#M��}�W�
YN� T��R�4'��2��d<�O8U;Fz��(=Pp���`L7��{K�{���[V��c<��/Z��L�s+{/v�_T)���T�X�Fl�:Y�z��sX��O*�ϼ��
�a/.s�R�@�����X��#�;)��<x���~��qg�"�:W�Ȱ��x���pB����� � 0��>%ӧc��������/�3���X���D^�-T�t��/�t���U���ڵ@��,gzj��W��O�unE��k2:9��(-y��p'�{͆�4J���_�^�Yn���I�vԳ�����Kb�)8�ȗٱ:�f"<+,d��Q���iL8AF֍˾c	x��O}�ʥ���j��K��o�Z�=�s#��]Ȫ�j��ײ?ǻ�o��������S�giy��T��.2lmfze��Q�涚��F+���X�.�*�|��T_G��X2[�n?��U�����F-�'�fz0���=Q ��ͦ�E�R9/���u�~&���2	*���q}���)���ȅ�sx
\ Ns�8vVU��6@��oa�]J邭l��)#�8�$�����.M9Jۅ�IH�o���\~��+/~��Y����ta�j���ҳTn'���8y�d�x�ռ����,uu`t��F��`�R��ZM[gSN*'al�#��]g���rj��ϕqS5~��MK�4;�:�;Px��Ƥ��L��z�L>)�����,���R7Ss}�z��R��͝B˒�6@wP�+��������0N�eb��#dK`�M��I}E��Lvgm����*Yz���?�Y�py�
�{ź�u��/O�*�ܢ>k��+�#�PA�wLyJ@5��,�|KWc5��V�-��{��z�LO�N�Ֆ��T=�{��l�����מ�\Y��K�O4>U�^�V�N����<^�-	,�������K&6�<2�+�zL�1\/jM~��ܩ��0��Y������y�������z�2y�����M�em�6�Z����GU1MK��U�Jx7m���u��3����@���`q�_}�BI
����U+p��Kb�R6rY��^#�v�͞��8`7��7�Կ�.����L�e�ߥ7��땂�n�f�UR��*s��pu?�ω������)����`T�WOS���}?QoөM�X��G�[GE�}o��VP)��RRQD	AZ:�c�!UDA@��D�T��n��y� ���]�Z�Z,�?��s�~���}�9wR�W�,�ˠۛ��&����G�"`�P� �>�Cw����>�[���^36���W����y����F�afRO�i����Xj�3I�o��lu����0��{`ڋ�zj��>�I�͑EN��+���7�&��Iw�Nɉ�B��~�o�|t�-_?戄�v��e��HH��d�e�U_����ӕwB�U�eH\�tU����D%v�0�EH������,��7=g_X}0�n�	[��C�B����S�'�{�2
A0"-h��]v�����m����E�6�Q���p�U��	���a���������r�1�ₖP�l�;�y���1~�bI�b��Z�X+��­~�M���%�t]��iv���v/���?|�ǲ�k��}0}�/����&O '�u�œ�<�l�#�R�G7����y���_Σ_����#�LCi��ܕe1K�Fl�5��3�*��L27���9QZ��+�L�RŁ�>��0�:�5��4��6-I^W2�I��"���+�/�1�%߿���c�G�������!�x���N�f��Q��ؙ��=��/<��b�-!5����.�p0�~p���*-�C��V`��8���`�C����Γ�������z��_�A������.��K���޳�V�w
�A��Vя*���p���2�s�%�6�a�ز�ӡw�~�WÄ�����?*5)�7<1?������d�P���x����dw(��T�� ��,X���$}���~�<�?�q=�7�Ӆ�/�IN��09,�_�?���߁�9�@�A����U�^�Zr�}����E��G1�n���@�'�;�8�o�!�����_ʃD�͋�@V]iߔ:DZ�-͆�v��b� L�8�$K��:j�;�Tȭ�R����9���?muH�
�"~�[��"4���Hq;�82J� p���ڶC���P�$�}k^'���ݓ��<5}"�W��W2��uf�^Uq��|�N��4=�&�gp��h�+Vo��V9�ٵ(�I���+�];�)��?]*���'�_\�Y�<�K[�}w�F���(��A����%�b�3���ʠ$��;�5�"_*A�(���Ε�[q-�%zS�Xe���P�o5}�o�7�crq�;��D���`���)Ef�o�kt�������:T��?���%6j��LP;u�WVB��q��K��9ȭ�Y��\?�J)M���c%�{�],"Pl�M��n,�%V'�z��OTU��_W�V���H�?rH��'
�T8#��3qq5T�{���ͫٞ"d�A�t�����*N�QS�Hc~�n��\���	� ���X=�1��xg}F����(��.��;;�DrXBz�u8@z(0<���̓:y�H���9Kf��>���~���r	h���[�*�~�����(�J��J戛�
��������&94����Nڪ}����Z.:��7x�pd�9:��zX��0dDKz���~C�˚�G��U�GȽo���Q�g�?v�&��[R�}x�����s���̵��c�/�{��������ݚ���1����v��_&"�|���+5I����_�-J��i����2��Ǉp�	V9}xO�5=�X5��pl�}"����|�)p�(f�{cX��/��5_|s����N�-�[�ooa�v:�;!�I{\#[�N�P��LoSm�0@/)/'�I	��Ȥ܏����:�*�Я�j��L}��@cM1��1��S�FK@/��&X@W,�œ#j�{.�"�$�Jɰ#r��omy�/���	+u׆�:ҋ�?��5蔿^S���
fJ���Ͼ��s��*Y�b�b�0m,T�S 5�����N
���@ORG�XO��9i���0���G΂*�7">,����֑v��������@�����r5����}��K���ͨ�?,��[Y�0|*�z��s��u��O�{H�^�e������ �5l"��\,���e-=qa�7��|�]��+����J��XL�0a����R�n���-�C(.2J)�� �7m������>c��g�^�'n�b"׼s�ɚ�c��3��7]P����=ZyȌ{F��/ɧu�S�We@ڝĚ�i52��'�=Q��maQߙ$x�Xo}_yK�dW�v|��o"ν�_���jE��ܠ�Q��GZ���:�pc�,�]����BRJ�I��B謄ui�s��F4�
v�������0z(�4��rқk��"�:A��I ��YI?�-8\��c����YH �27+yL�z�|�h��7��z�rD������_��S#Dɓ=�{�4Y�u��?������*�j����w A���w�
YG������g�¸8_؇��{+��P�w̐3�Iq��k'5��چ�W��CW^�1��rP2CP:�Q��X&:���Q�G�<U~I�_�K���������E�<pzs��S��<a�m6,&������U	������RM1�ֽ8a�8��q8^M�xh�D�CR5�$W~��W���?!��V���fy5*��)�~L�KuSRn�Oؓ����R��H�t~Z=AnW��)��S&i�d�6sk��h���1N�'#Vë��$�54��WƵ���(Т��M#����w�{��Ί�����Q�OO��z������e><���x(�H<0C^nT@�k>}��`�l�@�����V {tKQ �VQ`z�X缦��-ߢ�ҷ����M�>�p���:,HۻF�;y*�1<����B���޽��g"b>Y���0<?Y��{N��"�U��y������O�2M�Gu�V��)�����~}d����:[��7(?	�T��C��R��@�t���ڰ������}��́2�2�|�[_�+��~���5��8$��M謎��Qe�;�q����!��1b��r��O�F(}��}xeܟE�d�y���/QV�$6a�=�����_yxU���ە��bz�.G�tBi���
�W�XݴGߤ[�"`�EB8�~J��k�h�?��ghX�Q��!Ng�3��Nٱ��U.���U~Y�fO���з�:��h�!Xg�5_�1P�LA<�}�˩�!���F/�uL����`�gI���S��X�j�����5ź{ ��HC V�ȓ�ޥ�N�hǥ�h,� ���Y?�Ey�^������ۍ�	���lZ��u��S��zӛ^�8�v��:�_ƽ���@Sb�oNWRA����i|�蕎x�7����W��R2+�]����@����Bɶ���x1k�*�������x�:v���'�Nw{k��j����:���	�R~���K� ����1k0(z�!,D�)��w���<��"�7��J\׊�L~����s��B����@p��I��uL�63�T�h�+�"��h�I*'i���kR�s����xo�a�R`Q|�&���V�)�41��l>5A�yޜw/R:�F�1�S����N�vR�HC��t\��y��VE|[��
|t�����o[���#=�)PKh��,��&F���� �Μ�f��O��(9�'��[Oz�����5'��C3_�d��f��eߝJ%�����Z�Xެ˸�R�����@�x���Q���
0dkS`ޑf���ݾm�S�s��%A^g�c��2�1�meV�"�1�qf�v����j,�f���F�%b��)���8<���HS+CLVoC���_f�Mo�74���T$�ݛUxR����;$w�mx���\v��C��G�3?�v�#3��A. �x)t��_$Z�@3c0 ������9�������4���A'�@���܀dz��}�Y�7�*7��L7Ĩ"�;�e�J��F�:Eg�4�v���S+��Q�T,x��tv+��,��Ӊ��[�f���9\n��Ŗ�����DG��W�0����f��<���O:�F�J�p�$G0�:lM�	�M!��r�JzY��wAῥ���<�ڼ���"~A	��u:�VB*}���m껨�g�	/�Go4��ՉG��E\�?`��wd4V
�C)-���x�0I��K�eB<Ü�#���$��ώ������?_�w3`��Ƕ�(%�&���=K<��������h٫��/vew��_�u�|7���Yb��-�<|�a4�1�)�m�
��/���f�x[������p��
�ı�]������_�y��0�)3Jx���C?6�[��ޑ�q��
����n[Z��8��o��:�	��h����ȏ��K��ֶf,o�W����5J/��ٛ��u�?^���p!�,_-T�@~�N;/pK��>��^���l�BtP��[O1���(�v���,��9����y��9:1r2?=��[�)�'��+uٜ1��e�2C�{la�v�ߟX��Z�y-�YT�󺺇�[x�q�珠=���b����)�a6���j�R���
T��e��C�F5�9�Vw�NQ�ɪ���1.Ƽұ��Y�B<v>����q��S/�(�����}�~c&��;��"�O��� �g�~p�l��X�"y�Jü�^`�w��4�p��M�N���AI~��#s\ڸ"c�m~z����H���"E$e=w{����dQ���Cl��[qm��ݥXI��W�����X�VuI�X�V�u��m[�9�&�e��;W�?&>���h��?��_�*I�78=e>�|���s�	�B�8�9�� 1�g�s�u5�Aѡk���j�#��N	^��.���L�P����c�+�:#�6K,��^ޖڮO��"�"��[���1��Z6�s�0����"��:m'͇�j2�/68b����`�����](�9�#�#s4ڸ�UX'�����ee��qE~�zc��网cP-�����}>ъVn���N�`i41�n���.ԹXW�H�+��0>�O���_Iܵ��k�,�.���9cp�o�׬y�Z��V>]NlexE�
�X�}bW�O-YB���a�-�L�P���V�+�󭎩�!@�����=���U�����*�]`jM����ў
��wu��ĢR�H�j>���ʛ{3�Q��;֦�w�8Jo���:5�ɖ�k+�]�7��9�p��5��ŗyYQ��7�xe���J��*+��T�)�1���U�/G�{:iE�YJ/�3�V����e�5Y��C/a3"�,����%�ߐ3>m�BM�D�wD~��[�IG{��������[Smd~1��E��T�07/&�kS@#}��Ӄ����ra������f�O����i���K�AuÓ5�2�^�V>�����������F-�!�G6g�|������EG��jP�1mPTӞ�&,���y�{���94�Ԡ�jl?����s7�|�v'緈���掃4���9YRj��)��_E1�%���g��eTd65W��~�	W���]���͜窩>�rvg1˖�V��ޭ> @�]�B[]�Z�S3�O}�� -��7�\?��q�'G{4Ѝ ��y���>W��6��#ϧ�J�(��� �`�I��*h!P���ޙJ!��p��;)��Wk>��eЇ��W^�apn�l���D�{�ܜl\���fP_�h��Vsy-j��"X���_�L�Z� �h�9�{=VP��@T�2=�s��}��wz����Hg�������Z���2M�����9~�
��U����4�ߘH*0�'H���0����Y3ܴB1W�!��^�÷��砒�1����e�3ы-��OmS�C8�[�~�p-�Z�RR��wϡ�����rǡ%�G������|Z�=@>�e�����6��ig�0�[�c��RT��fw%���,P>�+����^[7V9�R��UIP`�}�x2�=Vbu\չ�}���*`���Xh�~`m�b,�
z���''.��>oh�;��Wϥf�XpzbR<�������\Z�D ��,��c�����l�3#��y�N�g5�.�y�vqE� XmT�M���9Yb�ƌ�;��h�HJ|E"�y�Z���$b[qr2z�5)�$`���x�wWk%����&���é�9 �0~�/}�(X+��gh#�P5��di�@����5�Oy��8����f����t���Rb�rKcѷ� ����>�hؤ���jȥA��+~U��<*g'Ն��0���*�6��NB�]���.���_,��5��}�� �'z�l_xu�ָ�-MY�������W��PH�h�����>5b?@sf��]����ٗ�i�J=AM�N�S�>n�$ӡ$�R(���ICąs`nwL����*��R�:c/^82�gaA��O��:MqM�eA�.$��J�P����0�K���z���`f�� r��˿d�u��	L��f� ^���a�e�#
�u%��>phYYBGU�&V�
ڢ�n?���u�nP)Ծ�yI��|}���Sy�l�)��8�u�毲/A�O!�Z_��-v�a�FI'�R�fڭ���:D�{>x���������Z3}д���3��wNab�i������_]ޅ-��:[ʮj�c!{��Q�L�A��zs�۷lc��D������Wա��(Ekh�p�Εq������:�� �N}�Ӽ�%GW��ق&��F�J`Z2��Y+s�pu��|�R����\i3�?jD�d%1s�&���O� �7ۨ�m'�U;�ټ���%�4�D���64ّ^�g�e�E���T�����{�L�^�3c��S������'Cb�2����d@���rdC�fx�����e,w�|	��Y���.Io��9Xp<)�lp��wb�r��n�Gl`�e<X��n)����-� 龜ص�w2�_qF����K4�7N�x�� ��b���8��8�C�'���H/�� =�m��k����Ӌ{s�? ��_��S��ヨ՞�í��n��TQZ��:�~�3��>c�=	H_����}o��q��҅*^+ٰ��U�ܱDl�y>��O��g��UlC1�ݱ��e�ZgM�&�H4L�x>�嚛5��ѿ��4�S`�����nl��S*��f�>}��wt��]���36�"#�yO�fsk!!�6ٗ�*��h�=9��[��-���^,7E�������������&�H�z�������,��|tr,2�]kŦ����R��<^���U�!�x@̲I��I�3YQ߬Q��5x�:ܰ�m����^HJΝU�ȘO�# �G);�]|����Z��L���-E[m�v�A��w	��v���EI&�V���^b�1��+)�g3)޷Um�Ӂ-=�E�+>3�.o��B�o-i�޵E!k吵� ż��y^da����~�2��f)���Z����������s�KN�e����w��s �Z�0�X,*(A@�y�����u��&�����)h���<�p���*�`u�,OM�X(�-�{���D8�D��jS#L2I�a��$�?r� ��Ԑv�l�H��;t�ϓ<�����^(l�;D�����@�2���Li�"���L��
*ڡ��~z"�)��b�Ƒ���%G��].P������&a<<kM���}�5cЎ}g�1��*�%6��>q#R�5��)���!�����E$t+i���k�p���7�o�}�*AݻQ'��'�G���K�j���9���Z3[̚I�X<�=�XA�����-�����_>���K�D�S����?��[�*�5s=����&~�IFW
��j�{��p��s�����Q ���Lγ\QrZ������{ Tb�K�y�ɴѡI.,��F�VxdbY%�t'�����]���ED ��1A~��)��QG���ϯ�-*�'��e%vJQ��ԡ�! 
�k�'x����/���š�FQ̒����(���3�@�?{��0���w�����Y���am[y(�8,w�#8�|�:Ȁ&�g�Vv���pr��i��5"�� ��_��P>W���&D���G���:��H:�|�/�4g:�/F)���K�v�����l֜ĭ!T
��W�9�٬�!>O.��|�;���׼Oz��.�d�"��:S�{�g+Tv�@{s�Sĭmoq�*U�\�� %)Gb���^?��e��!,g)��=��¯K�#�5T@P� %]�I��-پ3`3����2�|^��7�a�}��Jܡ�Y���!׀�دL�R���jU��lG��2�����N�F��u�|Ľ�@n|̷>V�y���L_��^Uh��X���j(��:�n}�d{�)��t<���l��H�#�g�z���ţ�V�{�B�/�Gݖ�j�uB���!�r���Xl��~�ֱ��=_ג�8V�,n���?���Xֳ�?MF'���t,�o��'80��-�u�1ԑ����SzF���1��M�2�;E��|�2�5B�2���L$�D��LOh��Wb���N��C!�b((�0>Oy�mH���5��L;���^D��_�����c���h�%���ύ���1h/򺇦���`zc�v�PѦ�{��Y2��C��|d�5e2�� M4h��!�fy3>�Mq���q�֑v�mގe�=��VV;/�sH�rBr����:�$!�Y��~�Z��h�TO(�1���a�wov��x������_����zI�	ڋ,�=-V�v]L�̄�zl(`��Y�C���Rנ��<��0qS�!-����db�r�ҫ�G���
Tc�Zׄ���j}�3�m@����vr�.buK�8� ��@���')�ΉI�C�_83��f�D�يN��|�E�
$T�;ʾ;�z��B��aߙF�R:Y�����F�2)x�|�I;�����kc^qR�$�~4x�ZKj���a�Q�6�����$�����x=���fT�'�����r�p 8�ݞ���X�'�At\|��$��7c��F��`�����lk8���6����U��v�&X��-q�4(k�I_&
�g?�~�W:��e�|��g���1?���^��"���]��9϶�U0>��ؾ���F�@v�k���Ov����^��b�Za�����@�e��ۑ�/��cD��G���%Yc��T#�h+�ͲA���3fƀ�ĉ%�@O2�f�(�U��v��ZL9��n��vNy�Bl@�M��I�ݽ�ޓIIr��3;��3��bD0HS��ط�N��6�(���P{�\������fj+}Le�զY�����k\�����uZ5'z4�<�[R`�o��t5�B����᳭��M�Y�>u$D+�L$�-*rB�G�O�H��	���o�O�#)R�Œ}����]m2Kf����
[�W�j�g�Vn)ۧ�8�\���؍
�(	�A��kٞQ8�  ��zt���%n�RQm^v�݄O��#QBd/��w�K��.�	�e9{��Dz<w�S<�%�_�Ր�	�v���C_�+/A�A��t����/���:NLd��+:���W�<S?NN|����ʄ�}c=��31vS-���[�e,��K֖�V6-��Jgk�b��sF0�x� hΓ��Uo�Ks���n�Bd�Ϲ%:6������W�Dh�Rx+�4X0\^�T<XL�l� u�}��[�,Y�E[r`(��,X:��N_�p���ɳ�a��O��ݻ>��.-����,o���L������Y��=.l�\��>^F}��D�tq�`���%$���ΩPQ��Z��]��E��1�"�7SDi|��UH�|�GY�:P(	�0N���\<�gip��t��b��E-`3��X���g*1G�I[�Ү�9'��E��!�pSX�j����f�h���`��� �������BU�tK�0-��`'{��G*�so03^�E���_�ꆮ��>ڕ�����TP��?q�?�X�JQ��F$a�h�#�Η��.����8F��_��3p����SK�Qʈ��C׭�my K�0I�=V�0��_�� �F�����Y N��Fov����K5����jF�U�m|,���	�pse�Ԩ?�z���Q���h���0����<,�|��=�4��mٳy��SG�����щi �`b�3s4�L�R����:��!k�2���)^D�si�%�]��9?%�u�?�@ �6���o�ke�����gȭ�6��h�?�0E���$E<`��0vy�B��] ��ۇ�M�>�Fh-※�Ia�a�zO�-8�(}���/����#�F�tS��X�)����J)A��y:p:� �1��)F5�7I���
���������g�ptíTE��{h'Í�T�Po����<O��{Y􉂑h�脳�dA���kZk�{��e}VH
|_^-�t�|uR,q>�(4{i�e�/�&�=K�:<�v�܅�U%N$^P��x�S1�F�Q4OvϻϨ!�Ake#��U�b�c���&�3+)�F����e;�s��j�[/ZX���ܵZU]�9żF�����nc�Ջ�'���[�J�g�&�"ZO��ٕV�WfτM�L�Z��uܮ�e_6�U2fqu}��Cz�&���K�hy�r���k�E�		ے5+Lh�MÑ��e��Y =�;�$��Q�?������?��|��49 \�m{V6ʮߨ���~$�%R�o�����o��Y��P���ӕ@����T��zC��f��Ͻ/����5-P��X�dBf~>��u�~w{\�s��P�½Rђ�yQ����IЩG�Y��|�7'����e3Ǟ4Q�T/
�ݚ��F����i �
0�ʣƳ�nqϑσ�d�1�%t��/���7��]��i8�b<�X+k �4z3g��'�Ɍ�E�����Y�Q�$�_]�`����2��꣹��˷�<���b a�mi��Qm'�A�����b��a�Ϗ��w�g��QqXr��T��s_ �����c/ஃ!=�W�ܼ\�"70vy��3���0�g�ٸ$���������d�Sϛ�:��-c�Uf�,���C�:����������|W;I��{�i{�������g�n���$~�/�G�?Eo�������ˮ��tg"@��^JHyEY�]���K�*��\��5����l�}[-�ϖ<l��J\>05�/�\k��-�����؝���䠐Թ�]�s�4�5Ņ�kh;=+¡��^�G��nu��N�D�T��~��~����7�z.�dF�qL&j���R�
��,T���k7�KG#:2@g���}&�z�5�x�U�m�i�	&`�l
����efa������+�]Y��1a�qiIv��^��7��u��$H�¡�xʁ7�;�8)E�V�E+������T�i�^�
βŻ^�&K�b&ׅ,r�$U_�`=�Q\�S��=KM�>6��h�EnB_����{ұ��W�uԡ��~��\��d�u%�Fz�v��v�HU���?�`��Y������ƁQP��F�������S��W��#qe����\/�����D}n�����*�37d7�ʕ�x�uj����ݤ|�P���O�ub_���[Q���r�n��Õ���]B��jH�;ގ>ߪ�L6�y��i}��s����f�G�Y��{���6�'�T�q��çvo ~��\:;y����cqEd��f�bz�B�p1��U���{Y�}YZ,)�M�H�y�7�cRo���sD�q��"��z�q�x�� ���?����h�V��{�]4���D*��G��������) ��e�Ϋ	�ل*ɒ����ؿ+Y�*L1�H�/�Q�O�9�_�@{U���1�޳\��&�����a����}0���� `������4�LX��#<E��EK{he��(-�S2Wj��B���[��>�#l���ߔJVB��ׅ]V�)�FD4j���ጾ���T��^��kw$d���4�:���_��	�83�4�5B<Z�up����,���1�9LQ(r�^MV�WY�)P�j���>b��;d�[���T65�� 2JV�K�3���8<��H]>���r�1/ ?n�O�ر.�����Nzt����R���O����W�Pn3S����m��]]���w�&��?���3*������%�5@��ñ�Pe�%���a���Z�5���� "��O����5C�E�B_a ��-rZ'��zMuH*Ƶ�=+�:K����j�y��g�o+��у=����iB��I�a@s����hϏ��Ƥ4��v<Ky��Θwۻ꧓��z�Fp����|Y>"������zn-Y���WIw��+�c�g\ _Ť�rLY�k{���8�B�����������d�z�Kc?�$��[R(Z��9R=zz��Bww6�B^l�\�!��U�� �;�y�O��w˛�?��<H�e�W�v8�K��BZ�A�wtf�;�@eem�����_�O9�.}01�*
�RÌ�,Wj�sJ�YJ��К���)��]L�~��]=�����w�}���Ώ�O�FW�}-���L�����\rpH�2��ր��+�O&����y7zC��> +ȃ���g�&��V�HV{������p�'yU'Q}�k�t�r?�}T7|[&���P��$�$��>L�'�<��
�(_��߯�S��KS_z)�ȇ�GP%FOߴ"�PF ��_�H3l�K��[�I��p{�%�n��.2��p�����١8� �t��E����c��"��ú(�mhW���--�TԎB�@j�����0�W1	�����x�:���n�-� 1�U͡��!�iYЮ$���ڱM0���X�����h=�
@�~�{�jf3}�w]"1��j�((��D�~#n^�R�|Oڠ�=C��9���Qꌕ0��+"�z����'3sd}��Xb���?����I9�u0[̸z ����d�����������өP�i��ux��R�a��O�[��
�񾺖�w*�z�
�?%v�qL�Ƕ�DP������B�,i��E���>����k�Y"q����?Kó4���E��5��I^�8���^��.2��ho<���ʞ|�Q�r8�hem�7M�zͬ��zl	u�������M�ǳ�u�d+V1���"*��ec�p$�����d8�348eyH��J����J5<ֽ�jrk����<�Ӓ�	��U[�t���M���Tߺɖ��A���k���(2�p(<�	@�ee��I�M+�����(���_F�,���0�p84з�R�e�t��)6a��3|yK�y�o�J����b��#����,����@�?�k�2lО�_�O���-��w�բ��u��$.-��⾓&a�o>C�/���>0��p�o� +*i�F��ҍ�"�0��B�~m��i���+*�#n<uc��&��ߗ�楒����//�A�wXR0��w��c܄��=�Q͇
�A�����A��w�XcX���+������������V<�n�t���7 ����X����s2=���BK�,y����h�l�0�sզW�����C��Ä���/�t�R��+0g��lar�gկ��eiӽ����O�q�mk���v�<�<�%�<�hy*-�}Mk��!�V��0�!��ֻ������k� A�eM����<�?�!�>3��Gg�.��X�&Pr���l�'l#U"vt�Ɍ���^(]�N�`)�����oJ_ѝ�����`�Bn��{�9j��c��T24x��L���-FX3R<���^�C_������0�Ӕ[���9�f�Gy�78�2��7�k!4�Z��酆�Gi�Ҝ�e?��/� ���޽����`��y�(-����h�ٟ)�L<��0��]�8]��f��U@�J��˦�~�d���o��ԟa��)T ���}a�w-��3���F��L�A��]�yo�Q~Cl���Y#��x��S��h�\%�ً;+r:,d4�*
X�tM�
�tP�Қ�\)�
��d��l���Ʀ���/k@a�<���p<_�l�NV�l�B[�
%J�����
�x�tz��n�o4�`��FϚX�)ZʶO�34֮��
=�~�e��t��r�u?.Epܣ�خ�P���U��Q��<�N���;w�\�ą��a������A�~�������NaTW���T��p�샳Ǡ�a��6�/�gI?(yf�yOV�ZD}����Cy��ݜ�I�����5n����e(����*V��ѹRɐ��2�rFg�s��ߤ?q)�	g�;���0�2a��&'�g>>�ٯ��S������C����(�;��=�ҡ����~./]�r/�'td(���^~�y�a��$6���!'���(x��n�8נ�������m���8␝"kje��Q�z�$���UR8��L?���}U;u�f�|��'�	5��,>ڒFy�L�{��hIJGu%E�06t	/Y'0�]���ݻ���D?Q�Lhu���=�g�8����<��ey4�3���B*����	��d.�[��������66l+��������-D��j�}���h;��X^��3㽹�#c$6����͔��U��<��~쵘~��ߤ��C���q�q��q
�l{�%l#�������猻�R؁�ԩb��~F�¨�A_@֯JOK�6"AZ�m���'�q��u�Ou��Z��?^�>�l�=(6���Ƚ��S�#/���F-�qȚ˰��/� ��w�,��{~�,�Z;�!�����(s�K�pv��� �?wI�A(n�1��8�M��d��\���P����v�W�G���0ه���jyz���fF{�I�M�dB�p�/�����"+2.��L�ͳ������{#����t�φ!<�cl�w�T0��X���h~��-��n\1nM �t�]p�~ YTgs�F�1�b�'������h�J�<za �0}�� �-dru}��e(Mw$l��M��F�:��$�|���qQ(�`�v�Fӏ�'L�O�ʣ�����p����mh)��ign��<�7��٫ҌF�Z_�4"Lb�,��
C�����u����3��9:t�Z�BP��h���Õ�2	�=h�Y^F�R��5�޲�	�ݫ�l�<���Mҥʻ���|�O��cK�!���sUe�T�_@w��
�H��G7c��V;r�7GЇ�PH����(��T�
��E#��"��7/4P)"��;E��q\H��z��K�e��u(���ti����Y��b��?�ɸ�c4g��\��o�ބ���L�n[4�<l���(=J��B��Z#���	��>�<[V���QY��9e�x\_�h
�_�8�ФzO�{�\>&k\7�ǥ�8/�FK�=:.�%�?0l����=N�/|��s�,��F���kZ���拫-���1�Ay��Y��ppT��G{��)ǭ�2O��w���'$�����D��u0�Ro��F���`���5{G�c���}�|�F��s"C��S���	#גs�R��Y��	9E䲲--��������38a�&����;�e �#���L݀�� ��j��n1�g�s~(`�
���L�>,��ѷ��E�'G��}��!��!`��;'o���_��]λ����Z嗵�5@��ſκ���.�NGLt�g��ͼT�`iݍ�=��xٚK�T�-�	d$�Rv��������`�W�J�����+R�~N��o�]n�<Z���g�����x����@�r�fe���̉I	ј�it�Y6���Y6_cOy��`��Q�����1�f���ᎏq/(��$1P>vc���O�����C��p�.Ӱ4���Pŀ ����"�#�in���F<�ү<����H�m�����}\�������
߅�H��Wq��kx�N�3O�t�i��6<��7���r���/O� ��5H����D������vS��M�Iq�y��P���l�9d�����p���,)�Xޤ�ﱡ�s��c<�I�Po)]Pk���
L�J��{�^t�y7*Yv�#u/��(��_|U�N!%�)KJ� ��g�UZ�{A�j��M12�_�8%�?f
��ԗ8S&c�D�i�@�*�Z��M��V�b��_'�7S����PY�3ӛ0�ú�I�;m���!�f
e��S���#�x5��%�~��P ��� +>&�oX�\_M�L4��{
	ޒ�Eܲ��� -���sV��V����N��j�g������[��X��s^���o���ը���{sw� �<��(ǉ<F5;" `c)V��`a-��pZ	C�fyWD=@װ���� U��9�&�x�OR�|��*�!~틄�s/�Ү���4�g3�
��9-ұ�F�-����h�B�v]�g�)�v��Ȫ���3���}��)�L�h�L��K��_g�{'�8w�{��q�}hR�?���Y�H�����VC����+M���I�vߡ;�ɭ�2l����|�rХ�|6T�J	���2�!i��w��������b�pqC�BU�2q�x�/����~2��N��Ca�3����S}�� q��{��,�����0f��B+1��Q�<��*�N f��1�U�yj��>���sl$z�@�*������i�h5�}��m��<�x�/u��h���)t��9����
�t���b���d�3EF9$S���c�ISxR4E�pH9n�����2ʑ��8r�PK\�����<�aխ[�E�9��� -|�1�&J��p_C5Lԟwh�ݙ�X����i���8axS^��k��]���`c#�Fp����'�VΈ&���>��b O������㱝��OdƎk�[l�����q��O���?駶�k��`�#H����p�o�������-�S��HDa�`=��S�����]�zw��l��;�p�JL���,Lwr�(���X������LЍ��O���3��ih�t��%BM���L����{"�ຍ�z
�~��OKʊ|5���+��Z��}��[�b������^�zz8��WREF=ػi�`}�q|]�|�����"�w�cO��E�o@�����7�c�S��}�73���_F0q����.�(��ge�}^�U�+|�Jn�v��rZ��!8ꟹ�Da�ގ��p�ΪD���;�I<������1�"��v�T�L���qM��.J����x���:<����^M�]�q���QaT�� �HA�n�HWi�T�5���
"MzJ�JP)�Ez�$@�B�=�2����޵d-��$'���{�'�	M�_XM(1>�� =T:�{3��m3������$���G�v������2E�����0c�-�[�C#�rӅ�R�_�[���/��I5٪�x!�d�&�Ύ)ah��M ;H�ޑ���Sۡ���/-\����߈�9�R�p}-R�1P2�[��%u�p�C�#�D��J~��B+��VMf�(�H��s|{0����/�.�m2W��3#f^H=?=qH0o<Ua��L��[������⻌��*�f}��<h��.����$n�M��5��T�QL��]�����}p��և�K<Z�ɼ�&��]�J�اT����^7���qz7Π��\]R�C��D�#K���p��I{���2H��<BG	߃��á)�:�����aIó��j���|�zh��ղ��R�v#���4��o���|�9��'�.�d�`�a��D�h�۩)�������[6�ߖ��}Ѯ�^�%]+�� �+O���=�����o�X��v��?|�ƪ�)�����!���S!�oFo+��&]u5_$>�׷�}ߓ��`o����i�^d��4y{ڜS��y�
$����G���ѓ&�C�Bg�3
e9�el�L�:_l��>����^�5�?��q��f� ��$�_a�ߞ��n�5)��~c�>�Ѫ'��U��J����ѥ;q􊐎;5vhR�J�by	�N�4(\X���`��I;�I�]@܂%Md���T�3�2jE�ij2����/��pV����!v)�O%"��eRA�É��e�iu0F���HW�U��M�7|Kܩ�G*���+�����5�����^:{	0NY�qC&
?qyo|���׈GWb�iAsz��=����臙�����T���F�i5�W!�y�mr�> ᤿sa�g�M�me�&��V���N�I��y���W�%�zG������?E3_k�ܙ�J-%�Җ[��[{��Y0T�E�2�3P�┌U�i�C�9�|, �;��_�n&}G��S|��`�w�i���p3ǭ)T7R��MUuB߃���c��6E�?H������B������_�x[h
�Ȑ)I�Ǩ
P��U��xz��s*|��ы���m:#>���/>���T���}5*ݧN�L\��|�C���%�0��))*/w�Yt����#���B��B�2�=u�G�v��T,�0�D����?bN�?��O�CG޸'?>
�˭�жh$[�Y�4:Zr�B��_`�EDi׹���ѝ����/_Np�LŊJ�M�h;�]�������o�Ve��6������H�'Ӿ�B�#����[zw��4�j|��У�� V�F�P`�H��R�i���s��lg�ZM6�0D5��Yp�0l�rv�咫z�0�E��W�?�Ƴ�V���8{\��n<歅u�.�<�]]w�H�)\�"���@U�?���!��x*1e34�K��V�R�z�-P�j��������Z�g�܇��}���52|P�3[Vj���G;6���h��[��{�-%%m���ΓIߕ?ԃ�fr�Bj�]���C��-���@��e��j���4d����b��߆RGK�_l�}��٠YN��^6����؍��I��'����������{.�F�g�3/��{;\��Ү�C��(�x+���N3��z�;��e� �x��^� �T�k5�~"b�D]i�'W�&�y�c��5��ª�O��[wbǆ��0+�kꝄ�F*"
,�W1ˠ�NxX��v��0��:*4#�UU1F~��<ǂh7=�A�zh1%"��3;���ݦ��i�#���W23���3�oy���d�f
��և
�E�F�
�/�/P��Q�����Ƀ(jBQ~�̔�`����h��f�2�gx�O\�s��Ja��RK��򊳒��	01Qѡ#�#u`b*db�+�_ͨ�t������C�
�H@fu�B����eYv�*s��kNn�t]������G(���%e�	���[owE��6R������R�`gz�9���ֹ�w8	Ɂoi�+�����?�#�p$H]w� s�{o:@-,�W V��W?��SF6��5c99���	���C2�	�@�>���2u5ժ�ϼɲ��8^�W�݈�On��=46TZ�Dg9)�Ε�Ӑ���#M���Z(���`5lTK˟���m������s�)�<��y#��.�:q�':kD'�ų�%�=p�:�B:]���������?�V���5�	4O�9W�a7�ﹹ9�e _���ɂ�����W���J��t˄8��b��n�=_���g4�yMK�W���DdZ�]��Qnntr�����A�T��f��	
�>��3Tga�hܷ
��o˴Z�� ���@�k���Ew�}|Z����l)��FJ��7H]�o�`�/�]zM���([zJ���d�����1\�E���7�H��DB�h���ϫ��{�֩ސ}�
����M	����Ѣ|�Й3h��NF��؛���YW���ɯg5���썢��
���V�Ţ|� |!�o�K��ؾL��ה�}�ᢵ_&�������dR��)��Y�h` ��f,�	w_t �T�J�PT�T&�b�I�g�X�,<����_+쌨�R(�5?a���o@v��
��u���r]�bG4���G"=F�]K[��28^r�k�X�V�bۭ��2���^�@��#�(J�eڀ%5��[�륍.ҩ��l^�!k_/[�^*Ȫ���x�1�݇��9�����?�!���20�͗�\�V�\�'m��WIώd�KS�I�uN?�x��u2�aXf[�FY�`���'�8ot,^BL��xɿ���\#~�K���n�Vj�E�!g��Ɠ�L�j�S�^E�^y������~k�.(C�y)���.��A">��ލ�(��,�3P�}�v���o@��W]��U9���ۦ�Uf�I�0[W�:--��W�9�g�>��!a(�<~���xR.K��M����2������ʇ�G}5���;����C{Z�~�G����t��%ԋ�
��rzߍ�t2�
��Q b��<�t��.ˍFD?�}�gzW�����٥��f��f^D��9R�:I���Jo�4h�n��'�S�,�����1�� ���$g�-��w"��`'Ҥ�ٸݝC�{�IUS=�\H�P.,4v���$�EE� �{�4E�������I�pL�����h��5��@?A�֋��xx�І�s���J������+!�o�t�K`+١ӣ�^t:�%$�3����^��z��Nwy3|:f�\Y�2�Yh�y2a�f؁�y���-Y��VJ��J�-����X}���EN]�g�[�7��K�>R������� ��Run��m�E�+�uN���7�	�24�zM�{Jڅ�<s�0Ev�-�V(G�4�t��`���n7K��HN=8^�S�ZE*����"��̕��}��N�O�A+B:֌nC�/�A	��������h_�Bgcц�E-͙�hkG*#/Ln�t=(��Q//:PnTN��S4���$Y��L1���y�.�0�_���X
ʞ��H�/��'�����v=�H���p|q�GP��jD��Z=��Ym;t���`~;��qH��z�ߗ-!?�Z1�0bS��2�J��v��9��>�P~�#�0�6�&�#��4jav��Yg�!k�7���$�t�Zy����羫��t�0!���M?�7���*��h����A����L|-�3&)�z���!Ǹ���֮�fC��AA�^A!,Y<В�"�R[h�6�M�� ���{�$�9cCy�f�߈�<x`ad�ꏞ���>f}e�;9��0�e<2�~w���K�>�V��L0�dC{u%�4���FU:2/����S��-�-*�i�]��<�u��[J���#Lj���aX���9q�(�
���`|�P�����ށ�ε�J���(I�e��Vg�ԞS9�x>�h�L�,3�u�|.�'�-'�vE�Á��<\uCU��<���%E8�4։��k9V4�,�3�.C��&�����Bڝ�S}���}�f���V�w/_^����q|��~�����Vm�o����8�Dp�z�o�x�:4u=umبb�߮Wq�� Uf#&�a9o۶�/��^JD�*;�ӽ���̈́ݰ�4�;�z�g��@@�;��"z�w�HK�@9����Ex�~9f��R.b�ژ'������ca����f���u�wN�BF����J|�J�w��M�+��#�Bh��/�4_��mESa�G� �_RT��T�"��&�e��|���F�I�����N����902S���[ƣ\��x� 2*��\�|�	/���n,�lkʰ;�S��e!=�m+��e떚��%���N�1�]����2@m��P����Ҩu�Y*�h����e^\��vL���r�b�Z�CA��j����{�/��7��4}Yar� GzASg�c3��^�Ϣ����Iq���
M����]�~90�4K<�yT�����4��nz���d��I��	���\���I�uӘ�߁���g��	3O\^�g֪�T��RB
�c:�A���`+`~��.�WɆ>���=pO�Z��k�gM�)0۸T
�WB�Hx��ݗ�1���M��AH˰!�xM{���]|o�*��Te��O����IlG�R��f	�l���)`̞k������KxY��SI���6��@~M��e��� �	�z㩘������7�_��1U��g ���8P�{IӽQh��.��%W=����A's�d`��_^�$�ἴ1��*�@�>Ogj��l��� ��yx�r�E5�z��3�����3.����������l�R�������4�m�n�{��tw�R��hb�i)�1-3/���(�H��λ��q�������U=�m���p�s�3���f;+[�_��qH��� n��q�:���e@��쎺 )GUj�՗tq���%>H��f9H�R��:7�����̌tNT�=�9���aer�IϿ�����Y>� �����o��@�4i.8/<�/�N%|�4����k�*�d!��[���\��d�V�>��~_MZ�i��{K�=��;9CD]�V]��M�|��N���,��`��9�\��rF��lk��
��BL��� #o����nW2D#v���#��Lm���Qf�ќt��qP��X��K\kQ� ��f�h�g8�|�@�]�W���v�q���|r�"��f烒
43�JGZ��َA�>�J��N�>oqWih�+s��Q���`uY��xg�(љE�� ��3l*f�9j�=G�J�w����66Yij�a�t���zs�dcl��;%���d��c':�G"�M��:(y�������͍/~�x�8f[SI@�[�8��دr��3O��Κ<0T��,�Gq7�)=�;�  ܩ`�V�X3��(իK
%��0f��2ᬾS�oP��>��^ܑ�U4,�	-ዼ�-��r�u]����b[[G/��6�b�E��MA�K$m�O؄�lc��)	�?J���X皀�BAO��E��o��;����b�Ө(ic�hW�3��u�_��4������<����w�Za�9C�}<��1COo��W�uZ�C_������cF?=�Z;OˤMwH`���EL1ui�"|Q M�Nк�Υr�i����S�C�A� 	�{o3�ݺ��bl����E�F��p~��h+��=���0��i&,�S37���X��mEN0���M:�b2�28@���� �չ���M!9�7��ϕ.W�;��#,-��et� ������h��\��يv��@H3�������ϱ�f.2��"3����)e�[W��D�H�`�<�e0���JDE^��`9ϱ�Jt$#%� �~��q��`�6&���=�k�V&G�tf�b� -�o�[Y@[�_^�}l�C�
i�-��}���X��g���gm�.�K m��l��]#k�W�.@�A�|�N������`��s>c��N�>�G��oF����@�� ��3٢�R�&E
b#?�[��[����� h,��f5G���� �9��y����9��b�SG���B�۸J1��Ui'�(׼=�ӥpn���r�Μ{M�y ����1��}�����4**bx8�*����%`��~hb`�Xz�� >^C��� ?����n^��@��~ ��ϭ���|�ix�~�����є�L�+Bjxa�b`ty�I�����萺�)yp5͋�����Z��̱k����_��}�T�'���5�3,ɤ���/I<c��|4��V�ݿ�ecK[ӈ����@�Te���L)�$)Zz;��D�:r���u)�ݾD�1�2)���}+��Dɴ e��{Q��e_�|m�̦|Nx8�U�r�B�5'E���˵��뎣0ѐ�o�Ѧ�#��p��m�vG���I���?MF� k��~��0���\s��4� �:"�-��i00� ������ ��vb^�����������(qW@�O�!��쪁v��m9\��S�]��e����0j�.�\ߤ�����֕� �zp</+�������$1�`���q�ps����+o��Z��߀	�c��@9#'c�8���i\ۮ 捾+$�P�-�Y��p~�E
�ݮ��mE�}�Z���.���J�ɀ�{IY���G&'������>{̕��@�{��P�Ց8����0[���0�C5��A�nd�Em����J�3ٞΧ�Hefui�)��K�˕� 򃛉�!���ݎ������88$��$P�������v�i(��$�r�(tE�d	�_��F�\����Phow.e)4�
���+����.����լ�2uvI�]F-' ]�����0��&�r�y'#������� E_��b����Ũ���� �� �ؠ[�����}�Ϙ�J�ĳ����]X���Į]%�@%=��w6�ץ�B~�Ěf6m�O�!�1��G"w�2���( �Q�6j�{���F�\ls|� K=�~f��T�s�;��27�(�uQm� ��l�]����}��q�@�h���\�$E�%�L�5G��)�&"��W���,l�5���pSz�(�252�@��]+�ny�!�Q��{֫�B�Xs��Ԗ�,��x[�x�hIk9�'0V��̬H�I[�&�I��.22g}
�ccL��M��l�/[a�0C�H��̎�}[W�����;-/��^�y��h�mM��$&�! #o�H���w��5�J����X_����!��ii�Lo4���¾<S���A��z:|�i�M3lz��49v�TL�J��{˝Q���?fS�b��Lإ��Q�h<���6�W��h�R<�+�%�\
ۉ�|5p�o����Ӈ7n���NsԨ6?؅z3N�J���<0�+���wVC����҇�©u%9Qs8׿�!I@�twl����5�Ԛ@����6���?��x�Ixcɓ)��n�Ɂ�����@���3h%���(^,�VL������x�UHl��PBkBƑ��a�sb�OM�P�5H�8=ݩ|Ҹ��R1V��\�S��6�Y����hP-�tѢ9|���X��I���C
4��I⯗	y�莩,��$���ߪ�&s�7�=�!OL��ݠ�v�S�Y�ň�.�f)��EL��,N�3��u���gij�����+�ʎp��yd�QU8�+��=����<��H�f'���@��6ZdT�^t¾z9P_RH�[*\�+CA]��9�>����x\jfwy%p����eͣy�UYam>���r'L|����Կ�,�d��7��d� ��X�G��;����t�V`'�����i��ȉ�Rb㘬ѫwo��!��h�wmT����R�$�@�+�6�������MŅ�؁3x���/����6SA��;vu����F)�p�Hb<�r��0�O~�S�d�U���H����J����{3�TfZ�i�
(l�Bv^w��2m�yۏ���� :׊�h�����d��bYLgju��k�6֜����G�U��L;:�W�M��}�*��FMlP�4*��U��eD��Ao��^��Vڱ��?�&?����!�����i����̙^�rY7d1$u���h�J	T��@-0�jn)�۪;�����V	�s�s )^?|+�h���N���W�Q�ٻ`�v�H��N�`T^�����v�i.�ÓJ��E�"~`:L�0��:��n�@��a&6�p�s�u��ڠ7�j�a��[��bGٺ�9���� ܈8���E�e����q�k��{�B�o P}�׾QgEN=c�"\⡺(��(3�V�b=���[�|+�8{p�h���m���*m�N��0w��0�UL=��f�^ی�9����!�9/9��m�'�[�p��u@���{]w�Uo���9��8�}��1�r��K�?�z�N�0b)��B+�z�M~����3k�{�z���tg��gŅT���T����L��HX�]���Đ�NJ0�<��Ɣ6��j4�	�ȋS���?�^��[.�]�g���� \�P%XX���V�	6�E0`pP��`���#�j
�L��4���x�Z���lgB�,9[l��w�f#xN��`LI��s��9�ڽ��'�C�����1d��y�m)gXr���ǫ.�I1���-��.�=�	���4�-E���:�+�,�<�V��Kq^�-��|��)~���=>E��~��P�.������M]�$�qd��ӯ�O�!w�_����E�"z������,���L��ϣ"h��w�J��ï��D)�dJ����e��uo|[<v֛>��0J�#���k�?dC�T��%wB��C/G1i�=w��3�d�;[�p��I���U78D�]�[�,�t��k���*M������ Fgef���c�1'�^]�����u����7��;w�˹�� ���'����BOy�������p���	�%)�w2�<t�#g*6�+�h�?>{냯ϸ�1�m��f�i�@cë���E������0v�6(ɔ�l4>U:Q���{�H���|!%Ui�����ks���n��4�_�L��'-�����B�QO�eۼEA��*kk�/<���yϽ�
�P\�
fm�yϋSr+�e%�z�rJ!���u�O2��QUP����{+��5x�-]�����~�'h`�2E�5T>��HX���Jq��3Tc@f}�\R���6�̒��`�E���J�`�w żyvA��H�\(.��zF��S\{����� ���fx߷��G���%�x�+�V�D�v��MX�� !y�2�$j��rr�[ )��SR�����6�2g��vC���[����B�+��]��C�'��:�����;��S��7� E�x+�oP��R�ߎjw_�Tќ����8��K�x+;J�r���lv�}_��!t�
6l����3Q�@"�v�Q�@���U�E��{<vr�˒���`?��/���_�m��`Ñ�FG���OIh����D�_ ��gP����[�<�4׽���^�]Ҹ	�žbd�:G�^z�m-m�.���������Ƣ|����%#r�ZCPq�	�X�@��Ѡ�������K���1v.�����!p��S)@�^w�����H��O6x����J�V���70�l)�R�[����cP� ư�,��&n����>�,܆���3�:O>����G�W��.5���(ے �,r�v�
NX�a�QZE|q�W��?�.Zڇnl���l�O�\e��SSe7� /�zGb���[�8��8�a)��	 �A��/�*N^�]}��zOiw!�<�W����$�#��|��]ï���'d���s�dN�Q4�v Wj��*yMM'<5\�6a� E�Gq���0���Ygl��<�©w�Z�°,�\.�BQ&������S�����5���7�/5h"��S�drO�=������7Վ=�z?yc�p,D�_õ~%�H�)�ͺ��U���B3� ��ƻ�^�P���{�P�Z����Rg}c��j"^�Op[%M-��L�v⮻�^+j�7.S�9Q�����}��ݏ�څĦ�.��@�e��g������I��VHг���Ȋ��rk����.�ԟ��b�jDN�ښ�3���X�?�&w���g�Db�Q��Lt�ju�2F������M���"����Ӛٻ	��@v�Al�2�"���7�+�*0Nq�=��-�f2�b�`���ޜ6H����
���'��]�u��O����\t��?YE!c.E�lIH�OM�{��X��Q!���%�p���l���ZS
���ۀF�9�WtlS̴�^��lL%)gp�kU����u���(�x���fYE��k��T�����l�A��r"���*~�'Csz}�)�<48g�ĥ�E!��g��E��e�����f�<�6�Vgژ�L��I���c�K�:W�YV���n�uo�������.���i,]�'��	�>ϥ����&��>0���"�b+Pp9=wt�F�`����-�k*��wQ��S+"sW?��ɥ���V�'yAqƊI��lM�,2���l����h�c���ʧ��p)�Ť��~��~�d��w`����)Ƴ������)~���5N?h6����o�Z=�a�WY��k����,��5�˰��ɑ�����gI=�vB];��<EARb��ō`��1�٭��
Y猨�-U�D��>��̜m� �M��ܾ<�r��J�����Bv4"��� �$���
a_A�̦̳S�L���HA��k�f�%�h���yn�T���G����^�chc��I0��SLc��6	��i�wz=�Zơ#��&-9JR��:@�V;��S$�?�0J1�0՞�u�i��WO�߇�E����hKjд�&w��e%Bf}����j�Sm[oyl#V�{�	�#�Q�;}��VC����I���<i	T�E%e��f[�����傑�J��(�U���)|ޘ
��{ "���n\����[�����!+a�b�:����RH2ä��7�]�� ��DX�V�&��Ɣ�:��e2�9���!��ȿ2��&y)v`D?�4�Z*��\ccm��B^@��x��!0�����я1BڌX���Ff�<Z�CcQ���gu�沬	���\uB������p�칑�����)�W�^�����W
�i�VO���U�ec�ٝI=��C��X��1Қ�G���J'a1����ŵ��A<~�$<L�ř��r�c����_�����t��QR�S֋���2-踹gaI�EH��&d�����l+���	߮���a��x���ͅ�๿�~:�G��_G�Ck.ZA_H�~��@��x��G�QY�Q<:L��΢�<�)�~�T�!ݼTu���:i�3���R�@�6�@�k)融�iX���ik���V0��=?,5в2\��Êc�הbV�H�=���zb�ϭm�A�奢��b��������8g�Ҹ�����)`=ᔢ&�Y��EM�w�6W�`i#�K��<�l��|�0.�����1>�	���J"��kTs��[p}�Z��T�B>n��}�.A�M�E��?!�4�)�H�^pߠ��d�N�H���H6�VM���#�gP����.E���ڝ�]ħ>E�u@�m��pX7D !n��3S�Z\#Ӹ+" *L�����s��\/VR��x� ��"�R�C����C%7@������gt��ʜ��Y�/�͟�%�����:I������ǀK#��&$�]����"�m{/Oas���Q��7!�l~�lKYԁ�_oOތt-�&dY�!و���L�^��8q6�Ǔ�+�/�1�V�FF$�������y^����:���E˚�[@k��� ��7�1 �r<�0�jl��AYqr���f�L�sP���UJɋ�R�)0G%I����3+�f0��� ִPI,2?x���O7�Ht�"ĬgQw�ND�n̖�O���1�X`���l���y�d�Im�)K3Ӷ�
1C����Ff�@Z���v����
Xyh��C5"S-���d����7�p�h�릵��C���Ӷ��`�u�B�r5-�Xͥ7��xN,1�Aӛk������o�5��j
w�E��nW�|f�:�$��%�C D+gF�ӻ�S�,�3��B��?0 ,����.�as�چ-���
9������.��d.�`�yBb�,����䳌B��z������Ŋ���FF�?��5&�N�Z�Ī;��EC���p&� !���D��IGM0��u�[�h!�q\��̀�T���[
�Y��W�܏ XZZzK'e~�jW���E��5i��j�Y����@
()&D���G�E����iӛ����BI���r@�j?KKԷ�k�Rz@vC�-�Ƶ�	��ǧk��Voy� �����y�� &8I"�qk�ύ�����z�q1!Lo�l[��l�'jƚԘJV|5�*ԙ�ؽ�䆱K��4��q3Ԑ�G�Ǳ��f�x�����F;�E��t�6.�u_PS܋rwe�c��rq�-���¼�����ߥ��:��&S��e���%ʴmt��X)6^�7�5q���S*�BW`��;2;7������ ��K���I�9����<��YKZM6�N(�$�l��-����G�d�Hvu��+a���(�G&u�9��^,B2��i�rM�JЅ_͋T�����5%K��D�����NH��{)DN<JY�J��� �]���$�Ku��vsa� �m���J��|Mdw��'v���u���iW����4�g������䞂�����l)݈k�I��pcC�6���&T�k�hWEV/�,�4���Ո(�Mm���~���\z�L�i_*%[�:�!����a�pg)�y/`�@���	�8~�&0�QiR�G�_$F-�xIFh2�����/��nY�x�Y'ֆe�_��������h���k�=�Ƒ���\����;���N�Bo`m��D�F���	<t�ݚ�5U�]${��m����kl0v;��v�O͸MΩ	�j��D���&�O����!�S�l��Y�Ԗ�q|�%���˄��VAw�KY<f2=9z�~n����z	!�"l����m�QQ��ޠ�+4ù.���_�L�Gٯ;�E4�;�`�9''A�"�$ݿ%[Ppi�QXx�s�U��	+˜S�GBr⺚��;��-Z�m��֊A�}���`���'���a��~]q6���Y�VRzI�b�&L�#g�K�� ��u˵�C�d�Ǥ?�ZK�mR�H7��Z\M��%�śQ?�H*�yJ�a��"&!"�g,�Z�ӓz2�g�������&3���GN���n�7�.�P��v%{�A���/u�kU���y9�� 76}>x�����	��]��v�ô�m�Ȇ,�ֶ5��6����fu����Gt�\ϋN%�B��b���{�j��ݼ_(,�)6����]�&��bp�},߅�N���#ؐ��������c����qQ+8���a��PŃ�s��؋��1ѩܤ,�Ȗ?A��#z����\�
�.[sg�Buv�������D˿},����c�5��f��1{M�0Y]`X�X1ݪ��*Ks�Bڧ�UD�/<�miHh#��*�T",��fjz��(4�70�|���TE�D�����m��h�}����F�,FcE%����F�/r� �e�Nd�h��0ę6�J���L�7���}��=�Cs*��,�C�F���G<��m�xh��%CE�|J`C�Uu���{�M���Q�m$?H������RSMp:--�3�b�¹A=7O}���'����������u��.
�,
]͵�'�̿{
�l_Q�b���f<TZ��4�y�]�F&���Ĵ�<eAQ��p�S2����r�k��q3�*��3[t���93ٗܖaxu}�y�$��>�c�y��ٍm��c(�^rxXC�ޛv�ʛP��k�`�0㚑�M(�Ƌ�����+�"�೵ZT^a8�쬏3l�x����aYb�*�����=���FD���"sB]��z��p�|�L+c���W�<��@GyJ�ڎe������OU��&QNƤ�Z>*��'����lp��ڃ�ԫ�(�LN2�g����L����_u���/������V[tbs-�����8tS&���&ͼ!����s���P�Q�i����������sǏZ�N����mep������m��͙,�K��﹪��($�2���^�}�ìbc����ɨ��\���G�e.�b�M��FZ�Sf�r������>��S�0ӯ";��M�v��ڀ#���#��;A)�/��6�]'�D����!�Qwv�����mYzn+Gs̝�J�u�,,Kpj�I��^9:(�[��`pin���{֑�*�nIC�5	n��1m��O��U���B���i�Z���ք(���Ֆ8��Q�ַ�!M��jV5�0�ײ}뇧iuŠ$+Նb��=��g�P�v9�'s���^��{�W�{�
�#�#�:Y��-]X������Es��u�e����I��(/�86��D��$�cRo��a�B�a�����D��7��1bի�aꏧ;�O�dSPU����6��6�������u�j���j����8W17���}���և�:n�R�fTG�d
�t�w��d�åֳ���ܱ
eڭ�.���r^�7���}ϊ�vb�!O|g�'�hJmլ�0M��:��,�}��QB�_�'m;�[�<8y�{=9�L��_�<�^4�Z�u�2�K1^Ȭ|�e"n^1�ΠOA?�Ro����n�WnFL�]>�bU�1�Ǻu͋��U/KRh��u+���(��l:����o̘�_9�����˛H�O�6��3K�0�M�tOi��n�PzJ�XhޜҀ�[���g�۫��=5u����c'�2}�:���f�x�;�7#\���}�j����zV6��n��y7�|��ʽIί���j��I��3b��U��z�:I�&�jO,!S�p�Q���n��ξ}h�=�>:3�,]�,IRYRA��<�usч�wC6�
#�
����
�W�����vi�����I#�Y��w�_�g����G�U�.�ޘF3{Z�^����Hߨ' Sw'm���Ч:�z9v0��>��ѥ�$��
=K�X7B[G��g�+6팷�����fw����L[>��2?��l9�B�^�����_?�i���������O������4M���'h���ץ���ژ�����8�������o?����E.�sџ��\��?��u�qj�����yY���=���_�����ϫ�W?�~^���y�����ϫ�W?�~^���y����ݫ�g���#��!����2Ō"��XrBvL�R��������z7�a�M{�C'9;?qg����y���V@�$t��<Ӿ��W�����Ϣ��j�Vz�>	i��y�鸖Ք���_1?��'k"���xc�۫�c.���qC��"��lj\��foN��>�ܯ���g��?_����^:�"�p�+k��=^c|�]�}�(�-��/[[(�gԢE��|��MȀ>WϿ���ԓ��Z��{�T�U���_"o�@�<j�7*���3��";������+�]f�p'�����7��0Ȭ}Gv�/��>j�Ӹ��N�����h2A5�f(��Ɔ*M��싽��F��^\9{d���ǎ<�S��G��h�ʌ��G{��e��d���9�,t�E�恻D�ŉ�4�B��%H!��hK��/�A�5�ۑ���ص!<�Բ#uO]����tt�h�ڷ��O��/+�h�Z�D"�q�4�� (��X���4v
����.D���i6�:�3{����?�����������@�_S���^���x� �B�m!@�e��xt���:k�����{7g�)A~�ٳ���7	<z��q:�?O��n\�eǎ�+����{(T��ީ/|�x���6t/,W���2�-�.��?����C��,��b��]��---r�hn�����蹑�hw<�5� �NЦ��v�W���!���f�NP��~@Ӝ�@�d�-������4Fkg�Ǐ�w�	ٗ�欣C��y1���#B�_w�h���O-�s�����3���3��P<ǃ���SU�B��h^o�ױ����B�\0�+�x"z�2��˗�hz� �Wn�&!�ko�st�T�ϓ+6���_��иi�6@K4WJ������N�����ʀ��˖����K �6����u���
��˗v��n}�L.����V-��B���4c7$׳�	�S�$Mss���_h~�w9�(X~�J�
�wo_�^:���v5��׉9����~��I炔���0p��#ݣl@2n±\���]�9j�r� `��΁^����v�D^^^�8}m7�pH��(mY���e��������I�srr*�oC���=+z�`^��h>���N��ksw�<�<��0z1���9���o{Fgc��F��^������2wss�s����G�Nt�,���{�N��Jhؕ*��!�����֓�k���SGg�ę$��tws��=�+.*�z�Ҟ���ny��E�wWrfff�i(o�eO��g��~w�ݺkԇQ�P�&�?0��p��.�l����w���Ԏ� 剿����u�S .�=V�W\H@����야]����(�u��^8��f���w�%��C�'
�m܀ҾVt7�n;���f0�����py�n_��+ X��A���ce:���s0 ���O�7Q��-�O?�ض�7�<6,چ��L�]t�h���	qC�nn>C�}u�ޫ%|���Z*���ސ��ׇ���S�Q���>3�AF;(�A1Vc5��(����3�m.[�YG��J���=���0E�|�� ���n^|K�r]{A��Ƌ/��������-,��*�$���YK%�8ǲ��hS t,��R�Z�:x�eb�@N�x�h��1�P`���;2zg������_�j5{��U1#��G	ͼ셯@q�|E[���ŵ�.D��9�'i@Z\BV	ьf�_���.���HÞҥ�4|�G���3@y񽯢o�8���պk�:/r�1��k�c�Pn���4-������ U�\����\'�K���{:b�I2W�I�p����ݹ��
t�Z��"�!���.�:u�!�k��s{�S�\�L�q�7`�GN'��v� �����׼nFiM�%�u$d�Tb��;��{��� U3V\B��AB}�?%�
�;z����Tj0d�K��d�U�l9S�L�X*+��z�4����{*�K�
�!���ج���t�-^<��=4>;��0�R�6>�� `�Zϵ����Зhܕ��\k	L���s�S�bF�QpppG�c��^�����f�+g�K����xUcOU��q͢6�t�����斁�
� ��+GUx������s���+�!I5;{�) ��W���F+>?���)��b�E�����.�Ɏ�G3:j�_��ɪ*�h е��Ȫ�D> y�w#/������z�6�ubIXԣ=3���bdx1ۅ@��Q�x9$iה!�مSuuzR���}�h����P�J8~�� X�!^�K���~�����):LG�|�W�/�IY\8����@�[���忴U�?ީ@�{cq�ͨ��*���)�^�yv��[����0ὠT��wC��@����D�!r��M�Rs;�%"�7�#��:XZ�CszΞ�� ����>2���H롍4m��y�� ���(U^�@����{�W� f�������Rjg�q�ǽ�����&��&�L~����+x�T:!�ڹ���(���O���|�Dc���2ю����:r�Hi��f	9�+h�\��s�`�{ (��� K:�h��h=��]QW��?FFcfgeݦB�w�4��C<�s��o��?(߀�N�נ���u4u}���V۪��VPQ�PG�BZQ	(���� dD�Rdoٴ�+��(�� ��^��B
2�)�Y"���G��O�ͽ��9�s�}�����Ԏ�:s|'�u |0�+/��P�@���b�t
�!a�O֞H��+y���kB��*�H���y��CCC��}
��h�#��NC5'	?t'b�<q��Tx���UM���K����!��5�J�QBg��2b���߉l���4�	��K����d��=i�B�脄�{wQ����U^)�6��:?�~P^�~��KM�18a1l<-c��s��B�֢M��`�O08�4k4%����'{�҃��<�&Ҁ��$�G�E����Bm��0M�byP�}�s���چ��5����/�Y���$�j��A-�c�87>�yP��ƉT0�W�b��ZJv�K�zB8ʽE-�̂�$����j	0}8yqee��<�S^�ްu��ya�k�v�� ��t��,��~9���љ����|�;Z�=7�{%�\��lI:�cVou�K�r�NP�z�:}!�8@lM�P�ߏ~�����TȓC�sK���(~�ܢ���zU�6C(������8ޫH�*�(=���hɿ�h9<\gH���&������S|lG"��_����z�,�׏/�{�f�`�Do�G��3��sIr8gOI�����LR?�C�XqvZZZ���|XY��a&��1�_㿑��c�G|v�0����̷^��! ��b�6P�LD��p{q��p�j���p���]v66��(�7��E�A������JRD]�>j*`��Z|Y���ZA�����:�e� ,[q��l����˗/�f*�H�������]{���D�۷og*��C-��Dݘ�
4��,����շbB�������1~JT!G�4��Ign�~(UsI*\�Z��>��sn���z�~p'��O�)mo��:b�w�Yd9K�A�uY�
������i�/c�/��P�z�s$�r���k�Vj%+yi�qC=A�V� ӕ	�˩��_K�mS<�n����	]L��_���r����Y�w=��s�^Z�'.���(ԣ�l��q$"�Z�ɞ��s]tՋ؊Y��,XK,��~��]������8P�&��g�*\�{�KjU�˚�E>4� ����/ 
��٭?�eu��h���/�����_9A�b>-|�;�zӥ��Q�b�)m���]��k��L�ݺu+��n�}�&�t�9�j楫O�2P�|~��
ग़��{�z��(��fR@���Ʊ6 7���Q�s�����v,�b���ήH��Gm�Rh�gP3�%�Ɨ@ܿ��Xp��^*fE��)�g�b�Og,BQ*c�V�a]V�}�ZT��
௮|���{aQ�H�7
s�Q�=�kOӏ���Nī�B�$2�e$O�"�#�J$�5�ķ.�SKR�J]�IQ�:�+m���ŽHZg��^��sS�ǗJ�>���*�F����Y�? ����)S�:����&E�����Vdu�-��u��`��8��7��DD݉��EB�,
Th`�~JK����#&�k���C�c��IE�Y^�S�n�Yȿ��1���"�B��ɉ�٭���R�{\�PW׮�@m��h�B��2������g<@6t����p>QVշ�k�{Rs�1;!ٲ힕Up�cL�����>�X_�#����m=�O��,�L��y?�qh�D ����x�Ȣ���J4^7���$2�3��y�� ��.Sf�s�*�^Ut��T�|	�$� Ԓ�H��Pd�U��k{{@�Yi6 �%��]q�Q�c���R��ϝ(#e撰������	���������ڴ���1z�r���=U��dH���ێ�>�	s�@���!��-���3+Zِ$�a��bQ���i�ROR50�]]],}���ϻ����ފ[��W%:��M��u�]��f@�~]V��m��#��;��y���J���i���mE�#65}�WQZ���!�F�JD52p�������*}���M�H��h6 f�u�rnh�K��Q�T���Ce��R��/gK� ����Ku���s��}��(�Q�˵�"O�t�O(o�&��;��E�] /;��ٝ�%A]�V(Z���ǇN���é��l$0|,��pL��GD��Jzv�FE]����YV��i5^UUe�N&��-o,^�߮��������?���O?��s��ӻ��o�0������[��m�O�*RRd�I����t��x��1�o'>�sݟ���[��ݚ'����V�8��������g�V�6`��n����-��;o��pa�2P������Vp�|��%T]��'���28��n׮�ݐN�U_��b�Ӹr��v1�o��|�-�k��Я�>T>��tP���� p�}�.*&�&�g�1��{�Z͖��v���e�}Z��-�P�إxz�z��<��;]b^�$'�^����l�AN��a\yx����߃�2;��{���A�Y�/.�2����cc��t�R˨��\�6��]�+�cnn��ś�`8T�l�|]wA(oԧM�6�����Y>���	P�(��#9��rVH.�5�a)+�u_������J�]-��]��Nŉ-�
��{��?�)ͦ����	W ���rC�E�Ы�x8�η���{��c�������m�]�֝���K�}�_\Т��{w�X���]@ለ�X'Eka��JVJ��#n����M݆��ޜ�*_􏀳#\�=�����7��,g���(����%�ٶv!�qOd��H��R5f�ϙ��Ǆu�0�z�)~T_@a�b�/�o����Y-3P,�u0g�΃ؔ�o��U���p�]�*ځ+�^��W�돤%'w�Zu�*��9�ϖ�%�m�=Au�y?ڐt������'W��Y��y��mQ�0�It\`GxǪCԄ5i��K�� ��G^��.�o"�n�Q�?9[UU;RkLYj��/�sK#[DmՂϖ���3s�;Kq�o���E�R��=��^�b[ب`�DTq����ڪjk�<��FUr�!\��#
dܳ�m� ����;���?O�6-4�����Sf�]�����T�s�Vm��^m���߼�߄4�`�B�q���w'���V���9P��!� �`>��M

;�(2x��`�b�'�Q+��>�АPᩖUɕ7��Hg�����F�����dCh�]K$�~H��c#�K�w4ݥF��7����'q�+��ii!����.P��}���;-xi���>}�t�i�x��8u�t��ԙE+Y�Z��EK�A�{��Q�gA����0{J�;���e��j�(h1�&�P��}�^�LcC�.�����	��G�v�F�Z�V;�Z�.�*��ҷ��-��Q�]�ioP���E^�cLvgSq�F��H�@���?��3��Ө���6��c�t���T�G�G��s�[�&�G8�zb	Lܠj�8��ꔀ��#%ȸ�6���º�11y����QN(x��ݼ�,P���2�5�b^�!��QG���\Ȳۉs�8+�y��O��m�7;oN���N>څ�?l��d^lb��\�GΉ�6�fbj:�B0^�t���Zr�)��z��X!Wp�nÕ+V��w�T�p	WUF����_�h�pP�㓑g������H~N]'�xT__�R�Ȼ����c�������Zń�ꪠ�"��8���`͖��k.��.�S�U���4�����75�<XJ0��ڂ��U���M��Q����u�{��$��$��q���*`hv]!@�&��'�}J�I6����!R�=��t��>>}+�=5D��6.�јӧO��u*T?�l��+����G��dge�>����T_�2�,H��ī�;��=��X�8@��@��n7h�M�f�vJTQhɯ�(����(5�)�N�x�g�N���]��8Mfˡ"z�k�|�pa6�G���ݶ5Q۬VZ��7)S#��ͳ��%�!�9���~��r���^�?�ª�F%�,Q��� ����HZ{���]�*�l�`�-��J4�f��y��0�j�L��˓D�hY��/�A��M����2��I�|߆Ϙ�B0�@�@eʡ�*�`32�T�uÖ_��9�#z@V��+��c��f�N*��fk�h�7rE^�yiMY���%{����vd׭����.�����/���5��>��!����27���ťK�"���è��S��ۘ=GP4���������WH��R�{2L����]��՘�gP�́c�ȕ��e�
�Tg�֨��7t63�(��{�����"by�W�7Ko1=L�hBcE8�B���WdT��6��f���Bmbх @	���|<۰�ɢ�`}��d yGҍ�+di�/��x������66A~��BL"�C9Q]�Eݾ���[�k�/Š�0�X�^�'�S5[��W06 �4�h�i�M�/��4�E
�F0W۲X"�j��"0+����q\�Q��"5��N�s�&��s��7�̝��r!��J6�6����:f9�.�T(�+�]�G�Q$�<0�kkk7e�]ܑ)w���I���eCǉ����S�t��%VU��վ[�]�o;��~MM�ac�@h���O�~?�$Q�*3Y��� T��/�If�ަ��Sk��& ?Nx[
UF�kJ1�t[Y�b4�ڏlɴ�����ɗ*��_II�g��k�Y�98.�`T���y�d�.Z�W��]!�y1=��{�<Nx�����eBN7 �|p���9/fϞmp�+d':�o�ْyQg�, d#L_ɼ�-�ȶ�F�_����WZ�b���M��w��6|��!��s�ہJ�Q7g ��Ǆ�����'OYʭ�L�	�Q�<a"�-I ��)[b������}�)zO�$���-�h�T�_�N{n(n*ޅq���@���Ċ�s	���"�;1�Gۚ&�p�Q{ ��:놀��LAM�~8 ���+���mJ��D>�\!_�?2\�Y�,�����:�0ݐ�q��1k�GƒH�����A�~�/���g�Y^����m1	U��T|1��r�d�y1{��h[�Y�P���ʷb���Ԣ&~�%���"��)�v�u%m�B�kC��ac3�S�e�3�g����t5�,'�r�$e����[�x�����4)�S���ԏ��dԈL�kz���HB�9fT�)[�lY}���=ᠼb9���k<u[{^^Z�62�5��ko��Ŭxf;�q�3���1F����TJ� =V�-�<�%M'���׽�=}\�_�H�n��������M9��g,JA��=I�⢒c�9ׯ��"�}N+��k�(s���E�ˆ.u���>����:n�q��ER�gk�+�'�@����8�c����Y�ui�� @������NTTT���VJ-p!��{�B7c��*�OeK�D8�o�fއH�P»>i��U$��N]$2��)�ϴwδ6\�@��/S�9���XY�����n��@!�ϻw?3�2����]뷳	g��%'��t�	�l���e�F�����6��b�����������:v�P���*$���455.p�YAH��YJ܋v�O/�^F��  *�D��W$&o�Ci�>W������G��� g��+�b�g�sR�q�+�;��d?rK8�#̑�6>�s��Դ?  ����)
͒z���
B���
���ԥ��b�$�}�����8����:�rEe����+o�@K��w�<e�1��w��F�H�[K]'���iklū�A�w�?�3��J�4�n��8�ɖ����V��mx�`�/uo�뱿<n`f{{{y����S��366�$�,c>%d����<�y�o:�I��̺N�e�چEdV���|u1K�{�33(�5\c^�%���S�\�[�;�nζ݆���U��b�^�� e*���V|vw����l1g}���E���v�eD�/(�f<�t����,��(�����g�����4�HkM(=�>Ė�^`���MU�dE)M�M�d'�)�Dlʮs�Ri?�*�o�<e��O��xrMnG��n���A���ӡ��ָ�M*`]w����u<o,�?e2#(H�ڿ��G�w"v%U>���ƶ�:O��5��΃�$Pt�1���q���$<lg2=ȆnRe������G+�C�
�%�d�B������6�`w��6+�$�5@�,!%�	��|�����dTw����<�L�P�������K���ҒK� �>�P%C�P�N���x���
K��7� 99��M�T�"�@�d�㤚�������,�ʎD�.u�UP��pߒ�zѬ2�ۙ��^�oN�3�r 磷nݚ��t�.��ؘ=vGTq|,d�<�_u�;cd[?�� YJ���7N����з�o�N��dk�ק��8l(9�S�Ʉb���n�0v%''����X�W��ُSy �Ѿ�ϋTZ��܇���q���6��u�,-����D��A�tU�o~�K���1a(\L:���*��n��Q��Aʫ:�3�����ġ���M��=�_+��B
�C6��X��V��J}��X�D�1����m�.��hZ&B�T��O����STY�d���G(o�� Ld}@{��n/�g��Qv����[˄]x'�{=�������Z��å��/����^�UdJҸ�����J���M�LQ����؍��ח������ �l(/�q|=�F0J���Nu�޽��j�$ֳLj%D�M��Q���c]{��h|/�'���Y�`!�����)�<����.��+1�ʰ�,�sf�@@a���g+r�Y��p����;�2�0����ƊɨĆ���	h`����D7r����B]}V5F��܂���x��̻p3j3����=
���Ҋ�)��S�>_���x�� ������7S�.]:@rA�*��^����ƴ���Tuuu�Ν;s����)Uk��l�A����0̀(5}h84���^��bɻj�d��u���DEiʧF��"��#�u�B�p0����,��p�c)p9��N~�zuvH��U^�iܭ�_��2(��<y�V��*u��{s.[�N�k����۷�$>/Po��m��
nE��G
��ћ�R5<�!��yͿN��1߼�;�sY��z$�o{F9X�up��J��^P����[,q�9�Q/}C��F$��U�.ģ"(�V�)oޣ����: ��ǅ�$��Bܷ煬���Z
3��U4�®\��x�&�]�jYG$|}��R�d<� CO�z�+�KP�BTyUT1͌�*��}�63�N�t�[(耱��s^I'5�=Æ��E���;�G�U!r���}�Cy| 	�Rj뷷Aq��o+jKp7�n����#G�MO��W�rr���yw>��g7��!G]��.hJkŶ_��e"NTu�KV302v��K7�8L`�M�r#���}�U�����Dj��[���p}��n�%[���Ե����tf�嘨� �u�T�d��T�
:���Kz�ަ�%)@=IH�e֥��m�+$����C��� fF&�\U��]���D��������^�wQ8MNWҏ
�����
�#�j����US�a�5����5�+���7�"Bh��>,!�@Ԥ �x�=��F����Y-|l�I����l�|^y�eQI"-�п_�Zm굛찗z,�A}}���ׯ�y!�ø�/�)yi��"�Z��ϰOJN�������R�,Wp�nWM�B+�'�`�߻E�i�/_�����7S�}���������?���L䋠l.��xN�P���&L�*�i�kթ�jX>�� ��?��|����q�0sQ���)��="[�[&?v12�]>{���6e㮹�ڰ�-ܰ,N����]��5���{{��΁��(�3�ȑN!{�����n�oaT!����Rp�l��ۦ��wf5�S!�NK�-��Z�|����m�ի��ғ���k��Ny��p������h��
^��l��Ч��8����*O�����-����:o<�L������W����v9ٔ��qz]�[��k?�	��+���P�� an(F�|�M��ꗓ����@L��Bסg5�Џ�Q����U��q��CNQgΘ6AY�h�Jw}no�f�|��#P����h�Mr��9���---�X-5|�K�����,0�Q�IgC&�}CI:��^O�����������x`�*��w,����kQ���+����o���;R��tr�=�$0}�
8�?��4���"�PKWB�{�T��$���� ���t�Jcb�V�C7����Z��ͨ�ZNkO8�	�ޘb�_�)ڽ�Ly�Q
vQ{��բ�&���C�4�[��ǅߣ��zq]����(8�Tqϕo�0Νp�t��������7�%Ӭ�|��:���IϦ����z�yP��yGv]�ɻQ��V�,�5������z���~���_�����}��m��H�%����:C8��z/_8\��t
(l<��)͡pR�RB�Ƽb�k^���6a;�g"�1�SL�]���X��L{��~�e%L6�T�o�E!_�G�I6���@�.P!oF��%<���i�7�CX�A���e����=T����
�j1�Ğ��W���������_p��Ř�;44T>�ب$�.�z�C���N����N�t���%ʽ��XQ��F�/ch���F���bz�U��yp���#����?����m�Z�Z^#V8߽Y]Scx��a[(^�ٓ��u���M*�tom+++5�F��S�5��o�S�^A�bh4�[��}�a����I߯k�>������Ǐ�ƻ�&d[��m9������%�	����d7�&'�Ȝ��E5O\�K�?c�w�xDl�'����o��k��%����.��9];>=��z�jӓ�x;|<���>n��Q���w�6;�KᗟL_�D���������Տ?���b����MI�V��}��g�4prCo���~zqq\y�]�>^�q�~���P&u��yς��֮'W��Hk=�S�c��Q�hr"/-ʂߠ�v��`(�5=%5:�{o���?d�ip����+:��а]�
=��]M9۹�d�(�� ^6��׮]�~:��o;���1&�b^!��W�A�Z6��kM2\�G�5[ʄ�{�V���5u�c�i�'�ne5��'^�� ��"�8Ա\p	uwC��V���Nߑo�=��b�X������	�B�&������q{ł��:j���*�3U-���7�ݖҗ�lM�[�r��8jkR����$.y����)�-�5 ��E͠.>07��dw5O|��%�Kq^!cP�<ǒ@����h�J��������*b���\�꾑�;HS���K��0��K6F��Bq� ��{��������P5>�r�A�]U2���?bl�.�b������%�J2H��=8&�Fo�����#��o~q����PwZ$�����v�q�B��o��+2��{,�IULy'˵a��)-w?!ݗ�&(��b]g�r�h���COf7��u�B9whSr�K��&
�āG�|��s8���'$�W�M���6�� ~^1�Q<f]i�w�P\x=V���#Vb�W��wdKf-���vttXI4��젶���U?4�<�p���B�Ԡ5�2UHiQX,��U^;eHw?)
)I���ZDf�]�6]�L�3=amL"X��n��Sb�L�W(�f6ct�R[V?	��	�:ګъl*J�toNx�F���]��鳐�b~���"�C���1:��הK��-^Ê��9�lb�.`63 ޙh�fwZ>����Q��2����|�&r ���fw]z���PC7��e��%�*�aR�����K0��PR�l������c��S�4��+$t�i��{�����ii�XܻE���\�;��V:��w��8ө&-�e3{Ɖ>�E���&𡜥���P�JĽO�=�q�˵�'U&G9���lw���óٮX۫���ϗ��
F��1�!�h˃H�Ȓ��\ID\	��/c�V�^�L�6[.є	V�!>anT[`����
[�*�sTvi��^د8��Q��q�#��g�T�=<���ᙟ�J��i�s�=��.fff���`B�Q��h�	��-̞��l�᫾�Ř�Ը̀	O!Z.QѢbg��Rg�,N�K��eq	��ϱ��U��~������v.��=���B��#�"E�̳����z�~'��$�1���K��JDi��W_�Ut��!KXխ���s���N_U��t�ҹ�ր�Y6��w�
.���mO��ɸ�!��kI�R�M{��P#�G
�H?�	��~�#a�&�W[�,lk�]3�Z��8�Dcj���BDQ�� MA��g�G�!��r��!u.ٝN1�ɥ�EQ�H�ݻ�������e5ڣ����g�N.�5�(����\�5���Ib34Jڵ���Sؕ�5}�P���م�d����Q'/h�s.+/O�ыS}!��R��j�����Mv;���m>q苢�y�a�ڏR�;����*�P��Z�w@*H�e��`�u���� ��Ѱ�7R���z�I��t��o$�.��r��C����v����Q��l��x���cǎ%��IJ`��1�CqS�u|��9uLv43?�w���x|��wX��D8���E���ܾm۶�h� 2�4D��S"��)�"�K����6�����x>)z�U��ʽt�1k�DԞ��ڳ�7}��sa䅸)ϯ�1�AP@=�
���Ak^=����Zo{*��G�leU�t8OQ�p����:��	���zf��N\�:��;���������ٓ^�A����r0T�n��T��C�^�0��Spir���%{5[\[�7<� o0�
ތ�5���R�־K��e��k��f����ɩ����+L�+Z����|����aެXc_���Ǵ�v�{�(�?���&'���kW���V�_��[���*���)��H�G�J�=/���	J���F�9,�1�[�nL��k�-�my!���ՖS;��	5~J�<ByP��L(̦8S�#�0���-����b��5����K�M�������Rw��5��Nÿŉ";���8h�3��*�+��fW꤀r��IPU\�r�{R��Rp-���ݚ�+��6*��<�%��7}�D*��G����X�0�KV�Ă ;�hCV܁�+��!,p�UU>�%op�^}u�� E�@z7a�Ժ��{\y$���>�ە����C�#G�*SRR"�Ʌ����n!�篢?���KC�_�]��ܨd�sNԻ��$:����+{�t%�{ʢN�3u�Ļ|���*N��\y�֘������K�y�fS;����`�~�w��З�x�ak���l	)|�=(�}x��yL�M��Y�I5
=���{孧�sv�ᆊQ� �����(>�����(�_�jD�!���52��S�u|/=�U��v�}�Z;������\�:ȥcg�V��� �Δ�%_�\������� �i���Ww�ګ3�5��ț��	Р2�����{����:YT�(�_���J	o"2��íڑ]l)
W�za{� :�PHΠ���s�5/���5���0���đ˩�cf�:��&�٭��U,*G*> �r}���P��CV̠QP0o����T�r'7��2�N!c�N(��._^�P�B�{���T�����L+/cם�Y�L��������Q�;G���F�9�"���L}����u��?M��^�	p�����M���G�G�$xpE�4ژ��0p��o���M����,wq��
�����ׯ_�K/~����\��
�U�&��&�cؒ�5���G���YM*u�}�U_*��K�����,D�#����4�ݱT�>��e�O�am�3�E�6ox襔;a�os"7�;�7�%�;���i���?`K�l(�c����z�t-�!��a���	ԌQ��m}�@�����A[j���E�l�����a������d���w4��h�_-�F/��]0[RC�U>E�{�߉���wL	/j��rK�޳�|r�Co���"�=o{�j�ʙ.��+��(\��݁6��.��%�R5G�($��;4��=_nrr#�f1���c��ΧJ:]L��cTMA^�p�p���9K�=.����S��4�J�l�]�v����+��wSݸ����Z��r_�9��<\���ˬ:EvH،57/Ѻ ۬�~��	�"%�-]�rd;Ⳕ^t�m8�4��9���G�}ZK���N��ZY�=%ō�9l�g�����>��J��S�4E���Sܔ1��|l��=>����0�*>?`иL�FH���t����c��*Z����P�Ol�̥���K��չ����n��V\y�&������̣��]oo����K�0kr��?<e>��YxM���dx+�CX�$�`TԻ��Jrp=�� U���n�P�X�x�l�0��\`b��U�D�#���ό�A.�ߌe0\X�Zy1ќ)��0��Q$L���w�$����OY��y�T��+ߎ��L.�hgʹ1_ߵ�[O�U	{��I��2y�}¢��v5["W���
��"���_��aDp彚-K�x�m�S�x���J%ͮ@�����%�r�u�6�^�K�u���!w���dC�P~U�����Iz�H��<f�qa�l3���\�Rzѹ���}�����-5[V���g�I�<Z�����؄���y��L��B�HW9�F��ֈ�6�*+f�;eq��oUEE�L⚟ӳm���z9Ӄ��D�����5�~z��5΍�u��)U[�R��
�C|L/����{<���PK>ڈ��m����֣n�Ѻ �\\k�������X=���CU߷#����@�@F��#�4Bx�az9p0���,_����������)�E�e�R��!C�!t��Ԡb��v�7�i�@F��"22�JN��v��/
�_(�����w9ò�/����ɬ������Ya�W�i��K�Z<��5a.SJGf�w^%�3a�;v	����`P�.cK��q_���%�8�ig�+�u�R�+�(26Y�%N��O�c�>��lieG����$F%K�v�԰߹s'�(8Z�NLW��)�g�� ���Y� �W~u��*��w{ ���PP����Ӈ����3>���r�l�UX���f����/����|M��Wrr�v�x��w'-����q���?ƒ���b��C�?7�t�W�B?��Ç��>���X	�3��wym�{�ҟG�܋��r.P� 2��〢'��'zBQ^�[Cq��,V�����^,�3�cH��Y�~_�z	���#�H!��&�H�Z�|l3:}�����U��Qq�>�+R�%0��V�x�O�(�~��*i@,���zy��"���%�X8�������h��\ya�]`�y%�k�lP�-�͑��:���i1��\g@�|C[�ʣNߦ�2eǄ�Dz�F�]vv�7�K/�p������a�"lQ�,�c�l�_�}�ї߀ĉ���Q(���j��]��xs�7?�5�
��]8��)}-�кn��Z���q��T�H� ��vL5���T��ܣ%s�OԽ�،W�O�˹\�ސ\�~O����9���y���o��F�p�pG�<�'��~l�y�EQ|S,<�}LOV��>|�+�E�F|�/�އs}69 ��C(܍��.
�����O �he5��nJ�̵	C�D)ަ�I�/`f�t?��w�M3q���Fe�kh0G�'�/�{�:�xM�W�o�K���H���,ta�?>H��&�|beU���8�u��g�S�
�s2������*�	T�G�-��D�)�X�x���|�Vԃ��+J������I���$X��;�
P�W+M��~�0ѹ��%�i<��u�]��e�'v͜�ξ����6���hk���~ژ=�`є�W�4t�@����������Ŭq7���C+V� E����q]�S�vO��W��IT���(���`�M���a¿���1���Ht��>R\�B�&�jP%R�b#^=��m��)Ӷ��qG�裱����Y��j�j��%�;K��k.��
���+�%d�d2��U-�@���	��f��,���j�����c��}Fs�q���>3���1����9�1M�V�+[Ҵ����*��
��Ԡ��7�^�!p�XX�&ܣ��Ɇ�{HE�}�kX5~Ёf�R&�sX��Q$��U�UP�� ]N��1��''����r���]��j��jN��
�����\v
�~�����n�
��(}��p#�P9rs��zcQ�>�JgL����E� ^����ü����� ����}�~D����v�l�|�Ԯ�v�'���N�;�Bx��ǫ2�����4��ܦ��T��&��dac9�}m�K�{�F+�`w�g�"L��w-z9DD��� ��ki��þ`�#m0I`�I��|�q���*G��LKk� �;=�fl��ڞ�Y��E�/h?�q��$9��S��K����hqW�v���l�/�|2�ri��6~�$����5��IK�*K�e\�������璓#�J�ٜ��̘r�#N������G�?�m��w�C̙���8�-����#!�:�ad܃���ӧ���;�Q�K�洽mʿGl�.��y�-�!8e�Q�� �p�fZ�O��}����0�z�^��P�Dq�
���/4wM>���0*hK�������.�����.mN�� ��hm���ҟ��k�K�GA�?(��l<�-�pʴLRE�r���MÄP?i*&�q���E,�MҞ�������5�9HP��P<G�Æ�(D�Sl�wSff�1,N�VO�w='g���� ^^|'�V֞x��y�C���9�VU5y}��';�X���a�J��C7<#/��P]�����H_�������f3Vs`���bʡ�h��ct�����:�+O①������dD濫L���0����|���ޭ�?����h��}| 3^�,2�M�:0f��-͕JHuK�A��k�z~ۇ��=�l��_�x�lԘ؃
;�>q���$$+t�YZY5�1ˏN `�����!�愨"$���[-F�VNڪB��S6�2�g��Jh.~��E�lk����{���i�ţoG�n&��~���n�;*l�\�9�M�bH�ю���U�����B�~z����=�NE�ǰ�/���jO�����?#NY�.]��ܘm�Հ�y��!�NX��8��$�1h~o��m��	߮�;�����u���X�����/�?^�v��L���e�Vf�H-]V��.���3su�Vtj�����2���{~������?~{�����_|�KzV��V�>s�m�ee>	^v���c��n.��ߏ��T=�v�knk�P�(��� ~��^��fS��Uq立�w|��ӑ]���ں���͏�]>খD䄗mC|�28��a��CZ�������/�������U�Y�Ϫ,�֞(��fVk;�|j�mc!і����^)(�i*�9����t=�Ws��!Gio��LII�(��d_�������rp��Gh�ϙ>�~�d4���zUdQ�����נ���]wtOjߟ�������0�TƥDGK��e�e0(/U�v�c�F\IttMϴc2�@]əE�.uq���F{�V���[g0���k9�@�M���{B�쬛~��L�řk]������F7�ÄB5�#�i�E���g�J�n?6S]�Mx�
C�E�Л���י=���f�X�D&*Й���Ꚛ��U�o�b��0yu�ʲ�\��UTT�f��t�f�����<{����1�m�D����0p���=N����@j��n �m����7�Um],�����w�.u�Q+�tX6o9nta"�d��rI�Z4�����\���,����2"}|���2=B������q���awV�=>�	n����r���˓��O@�-��gV*�:�������c%�o߾O�@W��MN1/��R݄�M�ԉ���������1����ze �g�����N���R ����0�"���<b:���������w_������cD�g�����}���$h��ߙv�/%>ř�%�%0h͂�a9F[f��Q+���5(�rZZZ��X�ƒP����C�
ʥ���wy�:��/e�,3��Fe���~��̣å��C7�S��V�Z~�d��vZ[x��(uM"Z�j������ $��9E�8W��qa�8�j�K]�݈}����������#��,�R�i��Fmt�HϨ7r;*@��4��-�k�]�,�Μ�7*�s�2u�S���r�ϛ����|��k/bE���s{U��+@���02$۶o�o�0{����L�2�=�ퟔg���X�u;��1��s����H�AT@a#@%���n���}��w��\V�M7��tC��2qɖa��ŉ����wE�2VH��i�'���ݘ��Բ��V�dե�,j��ӎ
��eb��ᗕZq�z�O 
L��0/�n�����'խ�hZ}�D��5��Q(�dPn�|i�TR�Ǌ؇����/���з�?��{�`�S�� :wxl�֓����87�D��T�_"����f�};�x�\�F)�hխcN�QeZ�ʼ��� U+����4�8T.C����;`��&������:t�`���!��[i����8O�R	>L�4���ΝC?���
�q�$��Nh $q2��tl<�ZDC�%��^��Npsr��HVK0n�1_W�_�	��4B��p�f��U�3]�=~��핽w"lg3��=��t�G4�J�`�?�c#��#�Ba7�Aҋ��u����n�r/�����`�6n�Xr	�
����g�W!#�.�.S��:s�<ح� s�3\v�d4{pՔϣ�NNN5��6��M�͏�Q�'������X��p�����S���+vM����3�%��(�^�m"'���*uC[~��y�9����E�dj�q�4�ٍ���r֜�0+�N.�h��兗��g��R2�����x�B�����W�O�N@���6��
Nt�����95��c��-��JF���9ȃ�K���P�y���:�>ʑ&z[P皟��߹��.ch5��R��酯l�v@��˟\g�<!t� o�`�G�.�%oRg�u�ԾlVK#Dw�W�ð������@�˺���K���#����s�D���U31SLe<4�TExE�u�ԫ��Zt�<<z�V���q$�<�R9bQ��@�@���Fm��BZ��n@iAJ��jp�Wto���6���VE�I�,�؈�cޓX�OW=D�����+���$x)���fy�y�b�a�
�;���IU�Cϣ�d�Ӻ8QPȍ1=�y�pa������zGN
�3�a���}~�L�ޘ�8�6)�u�N����R�\�v�֟y'P�e)��!ޟp &c]����� ���Zv@|���z�J����V��,Ѱ�z;([��:�4�7�~�ŉ���#@<v���	D�ƣ����|��Am��cr�A&~�ώg���yV���ͤ�P��d�P�oV(�Qv�7~�	p`�j����~�nH�����#>y�|�	��F�K]�;ɭ���"U&��h+�(������N�&��O�c.x&3��������7�t�BV�Z^���K�*X��'_)M���5��S����\ �b��+�l��&����E��[2�	�D����	��{č����������F|��0�?R9��~�`g���2�����x��) ��2P�h��$���1r�PX�f����?__�u��`��>�Њ�Oޛ�K���ֶ���Yih�9�}�o�хGG4[�P��2��~�/'�\|����Ka�R�������]��UUU��~���3�X�8;�1�^�(f�q���K����ւ��fc�}����t�A%�����p>����i�S�Oz�MR-~�٘ġ;B�h�������P��K4竇n��ރ9[�3>�t�X���vk���. ���� /}��
PoB�D�0�9���^=�e�`��9X�,�;6��mx��v�����%3׼�Z^��� �ܢ�u?|�|?�i��RSS�/�i��Q'e\ڿk�����)�{4!#�]�i_���.��:���a���{?���=�"�#KN� ,K�0�^�'w���P��;�-�[���)�C8����yv����vu�����n9��-�v6O	� 7�M�*O:��*7f�Ƃ��#�z�G��?㧏�p+'$����L�_�9n4 �h<�?��xAg�0�<ί�0g
�����5�r]V�� ī����� b'�L�
u�>��B���G��Ї\t�z�|����y,���UgMf#Ĭ�-�𽑁��t�릂�J�'������YL{��0|��s���9���'+��v�CQ}�Y����|�rPr��\�7��R�k@%Ow`��^h�� ���]��{�M�$�"��&_���'W>T]]���$
#5J������.u�$�vD�|d��
�qƑ�揭'�}gY��2�ָ��Y�;(�|��0��ɬ�*#ѱ�I�b��ə�����K��u��o�M��u{�ۨ+�@��-I@�ː0vFQQH��-zO���Z��0��Щ{S�)4�_��Ϳ�<���i�/����PK    {�X����<  �  /   images/bdd7c0cc-86d6-4eb9-abef-3fcf444ec41a.png�YeP^�'X��YX�C�$�������;X�ӥCJ�E�nI%�P����o��wg�93�g���͍��Q#1����H4ԕ���v����NI%��g=�M����z��~'C�Nzcw{��K,~'7o[��K~w/���2���4�
	��bz.k��wx;xq������[�����H�S�^��jz,��D���K��
9��+O��,T�"K��B��l�&�|?�u���YTT��1�2������3�a�!t��ư:��4��ޖ�[�\È��9�s(&�k��������]7]�ǃ�A�})$�%y�4�?u^d+�O�����k�Q�b��쫛�'�k0��b?�����ckJ�,�}��+�Kd5��Ҁ`͜�FJ h֊�d�OU�Yz$��D.��Ff�I�g+��\
1��{F�rV�7b��R����	��b~���&()�Rz�(����,��0��K�JQLD�9�R*H2��D��x�щR��㷸6ΞF>��U��a�q�Z�$Y~2�By�'6��ZQ2��`k$�bI�������p{]����1 v��X��f��2��7m�AKQt���L�;�{�Ե��h����czBSiH�D��!Ź��[La�����;˅x~\�%�f��T�ϖt��ߞ��ǩ��o���m��2l�f�:������>bE3^
�{�V��(a�r��^�.�L��)C�5{ǌ��!�?�W���ѝ>cl�4'�p���؊�g3+��G+`t��n����^V�L��4�}�DV����f�Pj ��޲dq�"m��BP^���[7�B7�\����7�:C6�=���\IIvZ�\����]�������
v��vG�,l���=?L
�0R=ƣ�S��8U���
�d� �?��>�[Nƻ�1���sLP@k����<�oD��ZY�U�\Q��q�\h�]� ���jnB�uk�I�ōre���<�ǀՉ(��^��/���3HԞ�b�M�-I��%+o�.���׍"K����hFt����}�a�����iiC�����7}O�6}�`���^st���Ƚ\�aB���TC 5a8Ԉ�,J�s#
������#�H�cS5G�|}�2����6�B9Z�I�&*֖_:��-i`�U=�1L����ӎW�o���p��<D0Va��qC���"X�_�/���7��dB�.���U"ST��u�(�;RQm�<4�E��c]��?Xfa 2��>�זY!����]��\d��d���9!ɐ�*�ѯ��o�9)�b��w�iF?a�
� ?������wY[X�߶:^OL8�-"+k�Fp?�f��M��]���v.Lع�O ����pL��g�,��&�L�릆�Qk#�C�]�g���*�_������N�F�G���i!U.�JlT��r��MDX	��J�L��p%����ƻa��k�>_� @��$��i�G-���_e|!o�Ш.�x�I{�XS�[5V�<0��`�X
�	,��RԝD`��6r"��Ya�[Ǌ&�+�����g��������^k��qBT~GG���Cޫ	�7T.�%=�Q�k�~z���_ǣ�u�*2�z��p(z������L�zkļ�Ŝ�#�����
e.6�$��O����ެ��	ZQ|��"Yz�	Qj�h�S������.�}3�����E�i�-��䲵��0MR;���<]Rd�d>Ɩ�c
�P�w�����ЂD}���{���zΒ��2�R7����;3��������w����9s���1����g���glS�87�*]�y�C�|6�Gg�4Ϊ�i�j?�3��i�9JuxT��f��� w7k)��YLY)�l�#1Y�D��u�-���*��>��!�@C��)�h��#��V"��?��Σ�d�?�r~R�S:��%�{m�F	};��Ě�c�c3z�}7ܽSa}��g5C���f�\Fr5�
�B?���(\v�7�/vI�⧥	3bb�^���������"&��,u���(�~���QD ���PJ�L�^� |䵖>L*� �'��Ԟ�URң�Gїv�Z����C�|2&.���ܮ:ۋ@�UX+�fG��Dn�m;,�oC�ݗ�{��/�p"��I��b��`�Ӯ�[�nXK�7a���!�WIې��j�*����eЦ����V�7��|i�ܴ�����фRO��/ţL��B� M(S���~��GVa>#u�����ӕ:DD��=�r�y� ���zi�D�� �Ò<� �J��it�e��т���+-L�:(�I"bZ8/�{�F`�i����1�j+�+!��qJO�B�ZM��ww/��-5¸��D�Ulv��z�2��!��P��G8��ZT���G��4����x2�#=�k4֍����O���V� ���pбe�ˎb�ǧW\�0s��<���{���Xa���:T�i����_�N5N�(��w�?=fd�w�Ƒ�ֿ]�|8�j�4F\'G߮�xً����a]0j�*�By�����@��1�L�����
?C~r�?���n����j�{�?��5�P�.G(]�8I�i�*2F5{�#��]�����l�X"ȓ�>So�&U��Jg7�^��GMd�`�@hhw�6�;[��1��YZ1)͍y���ǫ�q�l���S��-tMM����Ry�_�hf��Lf2�����4L����I2]�2�c6%�٤լ��s�ha�Iq�y�)%qP������ڿ)x��%�Զ11�x^��Da�t���`���x��H���;��c��20q?hv�4R��|�A��TK��4�"�����[������h|��hyg�߮P �J�ߞ�=,
낊$�\x����k�����W+Ԇ����(]�b@ER�J����������/�X,ү��b�	x���Mp�E��L��q �)TTlٿ�+�RC���a����"�v����.��66��϶b#���X��yNı��U�j4���ԥ�9���{I/S��Ola�A���}��Hԣ��Yg��5��p=8�)w�%�c�B�xyRLu��\5S�I=���BU��wْ�d���>�JC��_[s1�p�ˮ�(�Mkd�*k(x`0y���ϼce��"�JrU�_�6����X<��?"����ۄUD�Y��k� 	|a�A/�zЛ"����&��45p{�wo�7���˗�-�Y�63�n&�\�G)Ekq�#��b��S}i(`�\椨k�o��:/�'xL��.{���ǂ?���(i��p���R�$*�S�e��ͬ<���Е&9����d�*+Z�\���5�6)+��@�O�>���#�a�5(�}��?&���F����t�C4��p��Y�ݽ�0Dwdz۹��)KNؿ�&D����Y.����ʊⱢ���=J/�
��S����U[7���-p�AR��@�r,���t$MS�����XrZO�?(`)�֭R�H�i����]y20�EU"����=�Y�Xܭa�q&i",N�ɵ���j����]���������`YG��3��ڲ��*�ػ�y��~{M��@� ��:j?Ď,�3��7�頤~��1L��"���M��!�|'2�2����ʩT�۞meIR�xH����J�۶�E�Ĥe�Sj|j�݅������ �M�frP������n�U����<�C����]��@3z��Z=8Olֹn(�Z��Z����/i��C� �dݍ�N�>$��4�yp��o�rO^Yۈ�ԻB��Е�ސ�jFɉ��Ö�VYw�K���6����wYg<6���ɹ�d;~d���j�e�a��Ld`y8w�/��W/��Bl(h����ū�&�ATA(}�W܈��MIpT�>���m�uq� �l�^����R(]|��ݮ���i��Z��x�j6�j�L*�~��
�d�ꀯ�H��nq�G_2=_�螄�� ѕ7x.C��nyq$�R� �Uv�=eHF��cE�9)Q���m�M��&^^G���"�W#-5��x}=c��5X:7v$ԥ�>�,~Q4-#n�i۞�l��+X:TV<�ѣ8�xI��ε� ��Hr�3F�S��5���B������uQU6��Q����9"H�Zzk���l] ����4�K*n$��fg]:�%��ɹ�]X�Y�e�l^7}������hU�f�{�=�
M�r��^k,�^��5yn징k�Y������^���9�v�x7�~T�g����ʫ��n���p_�ʐyZ�� =��P{uz�6L�)�E8�����+� �^�h������j�UOs�R��t	�Y�\�J
����a� Gˊy��Q�xqq`I�~ 4&´���#�k>�M#6�Wb"w�����ڟ�VP�f+��h�1ֆ��������'Wy�6P�ei��Y0���w��L��@��ѱ0O��(z�p@U���`
��G~�Ӧ����pI�R
�f��F-��T�<�a:2%�^����4��
j�BP<�����=�&�W�������tn���y���1Ƌ�QF��_��.�8�s*_�՛�r��w�JG��Պ|g���+9ho�����9�ۙ��V@�fz��ȯ��u�}����Xq/k-���:q6M�H�欨�0R�T��q	�M�xf"���t��
.�B������/�*Q3����cẋ�dN���K�ǽS�bkFT^���"˼�����!kY]sQ�O����?s�r�U�G�a��2�^��ߥٹ���D�����f�p�ƌ7z^��$s$U���s�sfW�Y�+�X٫����?�SxN�;�� �%�L���yrny�e����`YNZ"�Ҁ�>�TEp��,��f�1N���DR�sD_~b�]�Q�|�`�6�+��bF���+kk���o�FV.��%9��7��}�G��n9q��@4.�}i�ܾ����z+l6E}��`_�,���V�q�o�up�e�� `�U<A��!?�P��tUe��u3?�q�"ʭJ®���@�TP2�s-p���,�O�VV�}�k�d��I;r�u���eOCơ���]�1��3rZ�l����q^$��Ǖ�r��D9�׭<EH��c�����'Mm�5^w��2�����}P#=l�1��I}�����꧵S����-M�d��͡�2�� øL:!�H!P���@ټ��ru}���:��S�s?��t�X��둧�bC=D|�5U��~��b����IH/��Ϋ>ݷ����Kc �J� �<�j⾔"�f~̑Iuҗ����C���"թL�C�_�LZ@�����זxf���(�В.�y;g&Д����P�2��H;�N��wQ].���t����J��XE܇���SRT�Z�j���ˮ�M!o!� cLS
U"~u�P�N�˻q��%o�~�"�a�����[�:�o��=�i=u��2�lHH'*�����͙��ï�w��H�3��c'Q7݉��������m��6���K��G{aK�(d��R�w�=��?�_�G���X��� ��Ǐ�&�' �5)����ߠ�œ�	�Q1u-\�5���x������������F���/hʤö��~ʉY��k��D�~� ��,F#N���Eĵ�����|X�=ԁ��'%ѝA�A��m�Ч��[�l^� ⷱ�����/��/K[��_I(��/���U)�Q���2w�y��mr�z�Jc��i�W�o����o��Z��fO�oi�6* ̳3Z�|��Ɩ��I�/���������4gt�S���~�aɒxn�6A����V��5S�5�=ZeC�1�W�S��ly�(���Z��K�r�N�C��2$��"}�g�F���N�u�hI��UZT�Ǘ���QJdgl�3���Z�l̐���&��U��?x��|���@��L+�U[�	P�i�U���Y�ݧKG��̡c��K���"��
�q�m'�T+���}����{��TY�3���/�z�Ș�>�E�"i.�z��w�����cW�1�o���ݴ�r�9�6�.?8���Me��*���?{A�E��c�bL
n��y��w�Jp���Խ�O��̷���X�����������#�T�5FP��b�����N�gO=3��+.�5��;�>��rɿ����=���'����H@��}N��U��3vտ�,�M�oTK�cX��VU�i����X�?0z@U!S+X���Зm���i k���O�Əzy6�x�",�XJWuU(�/S�����fM��F�������܌6�m�/(�n�Ѽ�ĉׂ�	�1��cf4D�#�6�lͫ���L���l�|E�
\R|�=珿_�Æ?1X�V(V�%7n�zح�*F�6@-�'�o��������*�����R�bϸ�j�Y/!ojݵgl�[�*E�
 ��Х0/��A���'Kd�+���^�,�_��0v����w�_�˝���~!�`�u~餍�s��x[�v{�Y�۟�8� �z�����MY�k��#Z�Wr�������N�vS�4���drI������Wh�,��ԋ�X�E�U3�8@������%2+�j���%������n��[)���+�Kǁ��3q �?��^֟u��N�S�N�Y�Ð�\�"��RQ׋�['��#�1��^�r���(�z�I�]i���4;2��ʙB��1p��[�Qno
 Q�+��u7Q|}g��lG� l�=������Ce?��޳@"_�L��X�l~~���Y5����?h�D���bD���U�a	��3��-��ۥld�gH��r�ޤč}�F���.�Q��E�i+$?��'r>��i�}�_׹b��Y�V�v�s����_�nk�J"#�N{h�{7}u!�����n��R3�s=|����/��s�˩@^7M����=��=x�級̢��a�{�.R'ٝ[ً!�!�L1�(�z��$z�����]����*�&��ŉ�T���1��N�3n���c����$�@��;�-��=�q�x�#�:^1�� �T�_�%`o}��?�����&2�}��:�5=����:4?�&���Z�&����:S�,2-d ��퓼Ɋ��р�JU���[!���{�'�gM��2��Z�}Kr���9��]�P�9��Ac���P�S��#�u�n^��sN*���à^���7�	ߕ�p>�l}�ӂ���Z'R�y��E�e�/'b�%@��3��Z���
��.����V�A�H�K-O����Õ�n]�it����6 ʆ�7Bo�'� �5H�vl�K�F��=Ԍn �F�c�i���̎~\���3�/"Z-���8��3p�z�}(�L�"|tYz~����?Kj`g�ע�		�
�x{��;s�$u9�+�Ĝ��|���}�]�
���׵X14�9�KO�E��=��?w���p�9�{i�ks���oip���Ww\�\��{�"XA=-c�b>����ǈi�����f�ǜ0:���sh�;����QC|+�U ���B��	��O���H\a'�N9%�[��c`n�c�N�rn�����۞��:�f�h�n�[vZ�_�)r�ۚ/1����S�í*	���W���hp͕�?�z­�����8ڸlx��d�i�:��/���zE���PK    {�X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK    {�XXs�銙 � /   images/cf59327f-2b20-4f20-97ad-1ec426c5b43a.pngl�T�m�6<Cw�t�Hݠ�(�(�H�H�HK�tww*#Hw)=4���>�s�k��Z,��c�s���M���2>5  �WUQ� З  �\,�'�~��oh.r�����/�E8�gl' �������.�C*WE}W]GKW����l]>�;}�u�l��� �
��=3�=<���1���/�U�Qq��hZ���DĊ2d��s>�u>EYẼ�SP����L�H:���pt� ;�y�o���P(C ���ȁ��e�$���)Й%vݚ �������f< �٭�=���:*�������0J��	���� Ԙ *@F��u��}$�)IzFf�Y�	��$��;��8d�+9������%F��-լ�u���{إk�o]s���W[�Zx��d�Y�9��$����ʹ��R����a�%燷[�2S������x�9�w;2z6,���2���� H���m�z�#�2"(���	�X�w� �/�q�լi<hk��.��\�X��$O�߉��s�g(�4'eh�j�w����Pښ�ᣔ��'�K�sI�NY7?ι�X^��2����D����/�<2��|�|���F��i�ŅƮ����5�H�Y+u�7	з\��NC�/�����dJ���:�^� z71���'"��gl�n$�n;{��h�t����u��va�"��bEie*�S�c�#m�t${F�滬�k�уQ�9��v��@�MW&~�[��l��Kl7��v�^ݧC�>-x5����n���,��XQ,�����Od:/z�γ��Z���Ol[��k�c�,.&�� �U��"���mކW�L�x0
�����w���MZ��P�0��-R) U2o�Ng�����dt40�R�r<�:��qݦ��L�,%]�+�ä��SvxA�mc��}��O�C�Φ�U�$�b>3�\t4 (gn���'`{�'7|�K��h
`h�F��[Q$*��4����@����d���55�y���=��$��n��NmgD�85f����!oc���_ز� 9L��)�)��1��G������ڈ�x�N��m�0e��/�-Ħ��T1ɝ˟p^"���� ²hHF.>M�<�n��C�#�d��YT������sۅSV�Zx�������fwD�ԼX�n������4z9���|�����e�2�hC�~L��c��Z�¢}�Ο�7o%�ð绡�p��}�v�=3�M���� v3o@�R��:�i�'^"������e)��u�����_�J2��R�d8��'�s:*�U[kj���_h>��gr����͛<K�>sN1	H�=0Y�r���{����$�^e`�E��"d4,�S	?��� x>{�_;�˚ě��������X�J��T2A�@�'�K�P$��Y���e�R�l�MR�$R�㺪B= ���o��EZ��8K��`�$�40���Cˊ@1\�Y�ӿ���'��-��e�Y{����Cv�:�m�V��o����mj��Ԑh>qz�'!j(�KO����gn4��JyC3�M��?��"��`��M}\����{�\{t\S.j�3Sst�߫��/�8T���3G����6�gj6����O�0�=�EЏP�A�v�#I�����>�����e�|��}�N	��¿���#��+ ��RY������/��W���K��\,����u�>�u�mUx�N��&�n���K�*ޙ{�L�e]]�˹���M���Jюt�+��^<y_e�<�[2{�8����@��AbZ�k٠<�:��V\����A������/�5EGg1c}	��=���%��~�ߍR��p�f/i~"�T�>�O��:�� tw��f�A/9�۽�d3K�X����mh
���_aߒ���;��^��˻1$~ZJ���}�rz�=p�e��w��/q��)�G��ބ��[�u��](�l��g��w^�8���tA��I
je���R,.t#�o�b+��ڔ�7����u��H<�I'�g�����(��Z~Nv�5��h]�1F�R�Ç�pw�$sC�6$K��q������t�ܭ��:Uq�-�AQ����?Ni5E��|�o�ڭ�5 �Ǩɿ睳���3ﵠ��� �ݓ��Aj�s�>��t�v;��\�����;�d��J֮�����P�8�-�{���Yz�OMGi��Z�������O�'�{�Ute�P@b��fO�C̷y�8c@���:�������M�G�X���6dտk\E�j����l�dʛʴ�/e@��0����o��8N��
���]x�)���5���!p~�i����-3���Р/8�r����>}m�#�4�1��A܍	;�0�-�M��a���%�� G�<����6��`ȏ5مt��u�WtF��{vhb�Ѝ10�h��	��A0� F,����4r�@;�Z��"ŎI�]�[e6�ޟ.�.�v�v����x}R<�_�)2���Ǒ~���ms!"�(>p��:g;������(��E�n*�����c�ͽ�k�mD���3Z��&��s^���p�e��d^�36,�sl[��S�8��U�+��_����EC������?r�٫�3�Lf��,m41��[��@��a��偳�/T�N���H0�F��v�6��8_�)"c�J+H�ǋ�;�u��@XƣF���������������i��$�ͧ.�<E��FbH��Y�t#�I��C����XJ�Ya�a60��p�:��޾�B���Ft�G�\��~_q��4�~�_Y�rt�/�D�8$��Y&d(�e��)z�po�sqA���/w"���/,�ܝrWC[X|8�����9p�LT�������O��7_�8��vd7�����~zN��+���E!�V�F��_���r��m�m{_&�z����˄�F�7;��+t��i��K��
�>`Xei^K������'N�Yh�W�D�&"��ٌ��yQ4%� �G$�K�?�yw}G9h	d1e�����-�<�:n0�x�;?���@������\ڶ�~B���l7���[A��ޫ'��g��љU~�B��㭊Ac~x����z���,ɼ	D�%m��廓��j"�x;X��|��4������]q�{fY'��;�,h��fe{�[��(!����L�b�=EϬ��δȏ��۫G@�Ԙ4�KJ=�9n<ߵ���hu\��uG;�d�/]�-�)W��NqB�E����d�]Ha#�?J��c�F��zZ ?�]���c,���VL"zlO�1*�&~mMݫK9Qw����S�K뎿�_I~r�g�c���m��)z��D�6֝������M�b�0���.�q�5�ܑ_��O5�>𩫅�'o"kE�]�q|�u׾����s��"3Wz���Dv�#N��G&qz/څ�U���P -+�k#���7=���Omݚ���%X�m̭��`�f[��̋�X�#|�!�������j�H:�j� ���$��9���2����l�8�#{VQ���$����I�Id:ȊI�.��)�����?����d30Naպ� �C�
���;:p,��׫�$`�13������SL��׈�j��[�Ƶ���wz���y/~X,�2v%Ae�[s�=�Bs�ܦQ�7�f�v�w�
���p=ח�N$b��+`ǹ��B2�;�،�ƛᲱ2S⋢����S�[�%���T�d����0�װo����>��}�b�w�t���4��F��kw��@�Ad�}�<��cmΖ�seʈ��O�w�\ľn����%eR��KLli� �5�C0	k5L�����I� �����A��i,茽YS|<�,L����e�hX��Tx�.�Rqd:��ғ��t��4�E����K
���ʀ���
b����AF.v��FV� ��Ewz}j�i��T�sz2Q��,c�QEY�e������lG�E}%���Oz� ��!���$_C���Q���ǃ�O��r?����1��6��W����u؇��L�����;u��zco69\h=���1)��}}�!�\׺m�28s�fVes����RNb+��>R����U�ǉ��'�4~ :*	*ޚ�+gϥ���S~v�$��-�Z?��O^�{�,��B]��@JC�����(�:�ެ�/V4-~�`I��9��c��
���ײ����X�k@� �m��q{&]�
�����Lp��_�KJ8�9�)tc�Ke�ےϔkl� �w&���d�UZ��I|��)H0Q��A��Zry>���ˊ˽�y1H���|�T�g�<����[�Xe�>mC���~�~ؕ��sz�������E+56Џ#\���L�X�>��d���o���/����E@Q��Wid�-� qt�n�y��+����X.mԚ��yҲ�d��l��B���]S"�&? }�䑑�M�޵�^��ؖwU�e,���h>b�?\�!���Ҍ��e���N1mqz^b�J��.��+D'j��(����n�(�O�[��;W�}����r��А�+����U��xI����������Q��9��[_�[�x����RUi���./��^��N��1=��~��;(݅Y�:Etl���(���� �̠1 �|$<80$K]j�ݰ6|`��x��L�)	o�td�<��P�{5OA�g��ݜ��72�,>�H�2Gz�x��k�2C+�/7�`��|�^p�fvڕ�l�3bVr���<]m�ø�W� ~GNV��z�#���"��LΜZ����1&gI��O���L~�j[��c.�e?�
��kMS��G�)�<e6နO�V�W���C�D��qL��E���ic��䯗����{�n>������˕H?�
��	�/�	�̽���3�i���:8{<��B[m9���=&YI�,�B��iz��<�=	���X�l����� �	�f8��1Dߔ�zޥ8M��T͔��tߤ������Kk�o��i��䳸���r���l?`� �5|��G�y#���*�i>ɒ�?}�'�N���2���֙���I����γ�兛dmB���ӟ�c��f-�<����'�[d�fzX��|B�����ϙw5�@v�c�~u�z�c��L�F�~�rd2\���d}��"�����9:}�I/w���)���L� �0@5c���z�.yϟ�c3od�N嫮��u�d=d6�囗��a�v����!�w�ܞ�)1s�u1�2�Ѥ��@�id�T�6�%i�Ef���ﴞ�U_d�k.��>Q$rz���gؽ��S�SQ���u��>��.6��1WvsKnsK9!��dZ�_��/e��$�wC�|��
�(��y�f�e9ܲ.:��l[�V��~�㸄V�IH�vvn��[~�/S���jyСl �jf��y�2>(�=�����&H\��%���{��t��	=�8��G֝�WP0?����/ ���o����d����ߋ9��\:��7�c�H^6x@�!;[?���v|�RC��1��R�& k�S�ud/�'3m����($U�L�'�Yh�����lCx�xƛ�֐���Q&\��U��TG�!-�5i���X��O��o<�B�u-�%�O:�C(�S��v�"{���͗���B݃W��W�)��?{���!��u5���>��7��dG]�r)b!+�AQ��>3q��VO����2!cPϕFv2�즪Ө(p���ӂ;v��/���S+�����J��?�0�Qj�u��xF�Q�R�c����HA:|�u�J�u����'Qe��7Ue�;"D�nL�f~4�M�5�1��l���2CX0��ݰb����E_�l��9��L��A˰��k�� �Ar����uzG�ӳ5��aQ 2��/t�j��5p�LF�i��YD�;�N
 �5chŏ�x>G'�hQ�9�L��uK�u���&���Y�t��[�f,J�M|�X��S�)9�;߄ĦD���C�Ԡ����a��y[�%��v���*�p)W�D�f�Q���a.XM4ף���{D�O@"V���Q;���������}��^��ɪO��hf)�gG��_��Nۋ�%��+��Tq�;?�c��'.��т~-��W��T�05)OpYփt�
L^��\�\mw�@���'k�Y���8�߄�Ғpy��A�R��*G�|M�h`�,�l5<����	�	h��/�Kr��"��A'�W������x���$N^,��0���؝�i����Xr�w=���*���Or[s��{�>;tI���E0��?�7��9j�R�p�)O=�f�U^�B&,��D°]w���O�tz�/�AoE�=<��d�%������+�Zд4����~�Q;I��
"�DM,�����أf������p�U�+�/\�L�^q���eGY���N��/qh�cKHwmC2%']�L�:0�Fe��f9��	 �&t���0o	�����)tZ�4�K�]�<���K�t���	c���߬�3F��K�(�<��%�bՖ�#J�齷%�@*���>�� ��#$�􆼝��&%���1���)&i��Z��`+w5��:ݍ���*f��ѿ�d�|?3,Ji�b���<^T����p�ņk��0�|����ۡ��܋S�W�>}>�y��+���v�#Ba�h�0��,�0�q��)�[�l���Dis$�)$>��7|�o*�X���?|9Gf?W]�ovmmJ��'ZW�HJ�bC�xٶ��\ \cNU<t�L���Z:ª���+��6k���v	�j�[����� K*5�`���	h�U7��S��]���1�o /���6kf��U9�J�;��Ӣ� o��`�>���4Ma�hd�`�_���2���\�Z�����ϸ���*^�]?lӎ��$�-�h��R�u�H�r����� ������bv�?�WU-�nV���d���w�T5�\JH���]XL徂����('��5ֈ�z���jjK�Y����Cr�����V1�rE����|)mR��4�m!	W����j{Z Bui(5w��lg���5뺂V~����8���k����#�ꜻUGe�U ��=}���+�U��q�`l��)��k���r�g4�ŕ��M��N�����5�E�1-�	%H0���'��Ƴ�A�{�9�C�����nf�,���cm2U��yI���c
.�T������7��F��R��3�u˪�d�h��ڋ�υ%Ju��}$S���D�	�&���,286X�5#G�q�>4)?{Q��.�ۋЎ8
�	>����:�] �̬�q�owZ�:�u��-�m݈8��� ������D�ñ��Ñz]i��l�"�[��?������k$��S׾���:�k"�
��w����& 	"T��
��۔�$T�h4/15�Z�Q���Fl�K��!An��ݷP~6���TPp�E9�W[ـVT�F��'|(��n��3ռL�e��}��짢�Ds��SK&��m��(�	t�j:ۦ"��.�m��aU�x�d�\��^.�����_�w�ӓ�dS�g/Cj`���_LB�:�m�F3�pd�M�C�����i��o>�Db��J��d�+B4N
��]&�;�ߠ�1C������z��.���l*3\���'8h�Ǒ)A���l)T��E0mT�᳑���;e���5:����N껫Wo�Yr}�����s9\6�>dj�T�xfd��^�=9��;��[��x��ONQ���E�3i�k�x�9�l���[e��O�4hl�e�_�QST�҄�����+�"�2n�j�F᎑�$��T��j���e�Q�"�H��wl����~so ���+����4׏�:���ʦ+�缬2k� d�M Bm�,�ΦMq��a��W��}B���BkM�;����;x��B_�㻢�>u��D�7�������ז�`Rk�H-)R��y�#N��	;sUFt�ө�6�$��Ƙ(X�葚�@����[����Y$m��Z�oK9?^�lgdOk� ǂ�
7?2StF4�[���n�pv����Ҷa�с�y�q#R+�)6�t+k>x�ѧ��ϰ�zQ���h8�55�sf1Qvk�v8�K�D�%�%!�.�G���|�HO,'����o��k�1��Ntdj�c�2@QY��S���^d��5�AH���a)W:/3�������P����=D����PK�G��CF��J�yk.��f��a�N�>�<H��(�z��8�!��M��vD���4Ř�Q6��Ӹ�	 (ԏ�Ea���������s	��"Ζ����!9N�q���)@���T����l]��i�;����u׹�K����ƺ]�>��7���e��^6�,ҷm]{
w��(�[���J2`���A>,����-%Rd}��.�G����QSP�R\�Ʀ}��E���y�)��)�ζ����֩����D~vO�[G�m7���<���a���H1���������q��������佌0�rdP�`m����c�e�O-����b��:�x�o]��C��ĻDs�$\Z+T��ij��;J=#F(����+%�(Mtej����o�U���e���"�%6q�C�F��q�L�__ѳ�y,[�o C~b�O��b��q��5̤��B���1:ZU�����|Ij�1&��xlj樝f��y\k��Ñ$�ʄ$��XQA}���گh��3��_����D��!h{h�zYO��l_����9P��m\�R0�F�y@�.!_.�k=]j��>8%�%�,]Ğ� ���+/Σ���̜�5����r��uL��r ��7Sc��:��0~T�p,L4�r�еSW�b�S�=#���Mô-��D�}�eؽy{@in����F������|��W��@TG�j�ͭ�9}܉���q�<�8����`�?X~-�q��U����%�D�39+�x��Rb��-^�:>�������;
"PყK!˻ER�5M)�r���l<�YD��w����p݁OZ).��A���S��s�D�Ɋ��ЁK!�␍*O-���s�{Ƚ����w�s0�s�kB�!&pfh����I'A%�1Z2�Or�\�]��j4�j�������-y%�%�o�K�b�H�}7\,��7����̡�M*F8������>�fM	y3]��'�zry9ǎ��sP���ђ�#�<��A���J�N��'Th����Wna������s���jѽ������9�))����l6�/!�m2D�mM��f�%F�d�#�O��ZoE�WQ;q\BP���u�t���)����l�z�7�ެ�)/-�s� �^�hH �����6�h�W�\Tյ~HS6��Y�ktl)��1l�z�������I�E�h~�5���殜;�;����i�衴3;�r�`υa�1 ��R���$A�[�%e}�fMQ)՝���hǉ۽��t��B���[�t�x/��
�����u�y��d� XU�n���H��S_,>jۥ|�?>@/������խg`�F�8�dy�2���_�bd��Q*2�xn:ۢ�d:���|�ޥ��L|��R1C9���9���;B}�l-.0�y������q�/d#�ц���4��o0���Tr��'B�����~2Nt�=1�[�a�Ù�bCx�[,>�M�lٱA67���,���oxĞ/����Db}��}�;����,}=u�_Q<`��|h���?����^r�3'���'����W��d#��o��
�}�`�,5D#��`�u����2�)9��SͧW��*���sJ�!�0sɈ���#Պ�1<6�]�
�I�p��0-EJ>kF=�f�;}��EaZK�����׀f�ʞ�8�_���'�hY��c.Ð��8�w���6~XUg��}(�I��#����r����c�fvM�Ͱi,�S��l�PH��������ټ�,�X�3|��D$��8��7��T�-��yBb�/"C�?�W�+f��T	�����T�0˻�^�1]S����`�Uf���l��a�w��+M�>!�g�e_nG���B*��H�G���d�>��/muZ�/�K��/
�̒�b O�y�[��,W�rkX��uT�B���S�.t�ĭ�3^5ݟB��@��J� S ���UM��7W������6�;aT?~@l8U�odK|�����! M/]�����^��u�~V��M�Gp%���}�����|�(�GTsJ��٩-�nV#����Ա����	�*�E�]Fng��"Œ�p�⮌Z0�C�V�qAj�Z|8d��viRSf�+;�r�������a�8i%��i)�qf&��H t�P����TL�$j��m�ޜ��w��Hf|Q46�V�f!5(뼕��c'nl�V���$^�`�^'�]���ۖ�X?'�W�E���q�[���-EtV�q	����J�H��/b�,v�p����3��=�!����hi�VU�4Ŵ��A��۹\��ɲ�F�E �+��06�C��#�H�1���up��p��L��|FaM�}�+�S�����,5Z�������="��ň�"��~K1[��9j�c䠥���i�Q�a��<_�7ft�8,�|�5~��њ���g�h�F>YvI���ѡ�왅�&����#�	�1j����J�xn��������-�=��J����=A�P�;�p�u)e�5Z�[�`���@�Ծ?��H��/��Fg�}��.�MM����{��?d����&�D;AF���o���^j_���e�$��Bs�띩
SA* /�e9b�J�P�����ԚY��iT�]n����|ᥦ$�d���?.�4\��M�PsE�
��E�(Q6���aE,�������u����`yd�
���e��7
�c�`��>a@x9$*L��_��w"��i�sؓ�஫�@�]��+�p�|A��'���Ռ�8aHfX`���|�H�W��/��n.{&cX��]�X�`�N\k��vB(K�D��I�ģ�n�"�zeͭ�A͖E�k9�We��d\���7�%uh`�dp`�}����k���Ԅ�X��/�U��~0�m�z�E���'��Lϛi.�O��S��t�w��J[=;ks#pSi1�����Q[�^! $8��������+�/*��ʼ�Vu��H��U�F�gK��軠5���5,]����}T:���+��%_���;��-�n~_���WO����^���j�1&R�G��#�.W	 W�YdQ��)�[�c��&��B��|M��*RO ���1��#��y��l�j�e;Y����%v�@������w��!�	�hc���d9�+m�-�TW�x�zkR���E΢j�5(U�5�|i�DOy³q��6�QID�v�6꒿�h��!�M�T�,���l����*��sd��_��X�bJ�ٝ�)�vQ���`cf�M�}���Q�/�d8�+)�/]���hfi�zox�Ϥ�c,ą�]L�`A��&���|��5i+m�_��o���א�qZ�������J�����>w�I6��ؐ
1t�=O�l���������ۀ��Q��3IJ#�ӽ��\k�b����rRϲF����fλviȌp��gt���I�.E���!^���"�zt
�����g�w��@G��v#6q�V>������Iߍ{^��Δ�<����h��yŠM!������(Q��E}("�z�����L��q�lJ��'"�v0"G���gm�+�pC���;�jTx��G�N���}l�Y��w��2�0�;��RF�����;f6�S�G|����ٗ
��^�� ?y�̈<&����r��y���e2�U$���U_���4�*�
,xH ')_��N-� dՀ^��vg�����!]���=66K���]���A��n|�9т�R��	=p�8'Ѳޫt��W��jp��u�d*g�Qh�M��*d��42�n����쓌���
-��ܿ4�>
�"OIȆujp��/�+���@�eJ$?.����u�n��J?P����z�͚΋�ss�o���T���ٞ���k�����ބH|���4Þ�h�,�#��ynL�q��A�`E�A䛵ܪDUשZ�8#Y�z��O9��+d�N}3:�R�p�|y�O��G[۶�����<�B^>:��dxБ3�����HW���S�<|�^���<�-F]�SϨm������"Co9�����]���g�'!C����X�����o��=�AQ&^A���8�ޥ��}�pN{��Vo�� r��@I�c!���br��䬛K�6�H�cb@�NS>�?cոx}}�уh�]Z�vGk����^�)lk6w���!�5��2Ic�99w�u�@rU+�g)�< � ����fGu$dH��_#�Մ[��OP	��`�g$���?�Na�r�ƿ	of_d�bVu �M�:�lK�aKbMy��V��0U$ ��f]�¢ϡ��p�@���6!�V�>/1 
O!;u����?�vV�A�P��']pz+th	��5o��B��l�P�ސ��58{�=醻[1��(}���!l�@����cY�3k�	Q*�KK?��1�d�&`�g���F8���)��?���KP1� {��MR2���bIz���/�"+�ُY�����^�M�[Fo�{�AQ6�(�oi���e��B?��o>I���*)��.H��aΑ{(�=$BP�8**
����޹�ɖ!ݯ5��@�9�>}���}��,�X�y#��.qz�̧�OE���jI^��}?���x�Jb�Q���@�Q��Ĥy����Luj��?����NG����\��r�$1E���"�O"4:�>���'�q���k��C��z*�l�2S�����>*Sǐ�i��-]o/��$NE3ػ��7Ф�+5��2l�x�jy��EF��4�;܂D~�vf�W���呺K�ٚ!P	���H�A��U}į��G0�K*=��}k���$�x��V�y�KN���=�)�����X���%�5���;f�c�o����J����¿��z�N�����k�g9H�!��R�/��KqU]�3b��w&��Z����Р���X��d˿���s��Qo8.h�9�o�֩��"�!�}����k�v5��1d|ωEW�W����E�	q�!����l�ŀ�=�_��u�%�":��dh�������B%������Ym��>�/I�̀n�ݔ���4i	���+0����D�'*@�����%���gL,m��8��
����d�����t�f����į�cüe��	U;�إۀǲ~A���v
Kjդ��ɕF�G�F7f�ҏ�	a9D&��W��͑��@�O��+.5N#-����n᡼#�gQι��;iR&����9+���*#00y[~7�����<�)^��k�ޮ������d	W#�Ҭ���*�>�\�n h5}����i��m�|���Aؠ?�F�G��� ;���8ݲn���-˥����,U�,��w�����dj9���aai�P�N�&��2MC�������,E�����NxlA��HH�>�5[[)pz��)����w��m���g�4���&���%����eŞ��g&-t��6���������"�P���Ba|�D�'7N*0Ա���/��}���"�:r�Zo����^�a�
�@�E.]���ہ�ޏ g�}��^�M�O�����˹k���8fi�ܲ�O�5kY
�э�/�Y��F?<;(�դs�!�J����'�/q�:c-�>�:[?i�6i˯v�8t>�'��gs���Dn� �&��s��ڐY�k�|	����5�I��9�ɶ.;��,Ňo�S:�5-�뗹8].�goO��,�����^�<�ey��ړ����~�]���eYh�t��n���hj���/_��ez�9!��s7�A3�μ��{\���4��g�7R�xU��6k��\��V _���,�4SP���`�yȒ�b�\T:�K�W<�nI�IHD�3Y~r����ca힋�}(����TV������t
���~�P�P}�u���oa�W�O�ϰ t�<|�����5%?�5������%���}�M�k=�P�����m�+2��������i"�^�./V�'���؛���o��;�_��4�H������f����:�1�["�k1��X�{�s]_
�e�ۧ;AL'm.�$LN�I�[Am.QBK,i���mwҬՐ}��9�����M^��ꓜ�(t���}l�3 D�A���� �i�Ub��j�����}������ĝ��-c ����p�N�D�<����3<Zj:~���sϏ��?���E6Ndڎf��N��x)OK��4����7�k�o,�f�ŇG��"�ӿ��$w��	u��0.���}�Ԁ�q�����F��'�N��@Eb:+���](�������+�h�o
Y��Y��9���is�h�5|������k��NtR���ᡫ���^p�ʖ�*g���r` Ï��l��Td�ڈ� �` ڳWI����9
�(e������_�%��β�i_�����l���ƙn)#���`���
�|�#�!Ig�5���N�e��ޘ��qM�N�p�=$F���_j��2o_�M�/p���y�SFi�wԈ���u�q�c�ј�A�p;ӀR�S2pl�+L%@�:��.f�l#�����鮀�( ��iC�-��}��B5S������1%�ʲ�[�t1�`}|��q�WI��Y-3n�oI�hڿG�m��$R�kʪF������>?;�w�����sx*���%�(�u'��I%���S�R_�B*����{��4O�%ݘFmo-K��?�&���?���\-��-j���;�)��q)2E
RPh$:���:�Az���>���M4]��#�3(!֛�a���L�ՔH�V/�lu��y��bn�1�l��sS��\|��ac�{����\��c��1�RΆSU�uS�_��8蓎��r�)�A~�.�{��<�tn�}8�M*v>�T���P��<D%��s���](�:��̍�W�궰'D��ʢ���v{��SGT�#��Sm�EC�p�2 ���|.�B�w�(��Բ�)Sa�툩1R�/j�kQ��NF5Q h-#.N���� ��UE�U/��Kc�A7N�Ys'�
Ǖ����>�A�?�C�J��(DpL}��uʭ�t�;C�=6f1ss���$r\���wZW���(裒C|!���zm�I��v�F��y�dK5a�tiC�� ��Y�ﻹ�	;�rj�#�2[Jf�a�#$�ȧC&z�����o%hొsq0�{��/T��'.���~D������J�A<��a���?}��{�������<쉂�Ee�`y�*��-�e[9�b/M���߼۩n
}\��a%��OD�借V-{Euh�.UI��
� �6�R�<9w������H8c�,f����ɡg�3âUS-'�ZhpD��N��b~��!|��'�UZ��b��NQ�*�Cs���ΰ&B�*�ks, ��%oo6����a��M�ڣ��r��qc'�lgCRT��K�Ñ�v�"��?��S�d��X
 0?=����%J�#�g��a�y���'�!4򌋏w�uK�#^w����?fVFl+�,��H�J�^��.;G\ۂ�~�n�%y��@�y+>K2��{�ZX��m��`:�[1����樦�V��S)��w�����t]?�G^l����~�NS��S��sM�a$G���F��푢�pF}`M���t�[�Nٱ��k�Ț?b���BK"_a���ڡ�����|�s#i`�&.no
�~�4� j��"]_.zI�]`}��|���2���a~�h]�z�A���c��W��8�	ׯ$��T�F&���L�� ��V(�q�Q��Ӡ�`�?�&���f	��(^_d/lXe$�~���#q��>�h-Rd�ޠ�Q�R��<��5A����NYc�Gx)���V�O@���A�w1T�Ǟ*����.������߱�i_?�-3T��PD_�NU�������V������AfL��H�v���Xib�5 ���h,fۣo3"��bzFz^Ѡm�`9�	�"��Zؖ:{-�o��������G��&�BU�TƱ��ܷ͠}Õ�������d:��/�*�\neW���eL^�ĭmh�Jq��/�s{D�Hiz��v*<A��_W%v �A���ϐ�B3�j&D���;V�y��7�A���)�?P���/��|NtX��6u����
6l#���(�:��g��qX���ͯ�T�]�5�d��ύAQ�\� �Z4,sm��=��Ab7��R��j%�1�J���/�1���mAX��z��k?���t�F%_�'6�W��8�"��w���O9���ޞ�e�v{�����au^*͢���&��f�K���?1ahs�����렠ka[v������GJ��������2["S�/S����ݫJ�[L�����d��T]�ȭ�WU�0j���0�f�Z�'�H�lnņ\�����V^/1y�U�r�� [�%K'A��C,<�伥4�ew�c�U�k��A�7q��Z��䯷���T�c�V�y�
��.�;�h��#�P�J��I�4�z�܁�� ����qQ}���0�t#!ݠ�t���H#�Hw��4�]�4Jw�4 � �����}��f�ٱֳ�z����l�[{p���lek�!�_8����ym���Bq���,�"��vr�M�Q�|�U���Od�h\ҧ��Ӣ�̳7�*5�;dP����:�v׹�|od�|n�ž�e$�~�"�1�qw���H��>��j�#��J�s�E'��~T%}H/���56�/�=��2�����wL�_'}墄��C�F�ۨ�I�@���[�w��q��Nb���[��麱s���H�z���p��/{��&��P�09��Nx?[���J�6�� )�$O��#K=�M�C3P�r/�n��:�ov7��cc�n��CD��u��v�0�^>)��gm�&Ŧ�=��0�/��u���4�7���^����#����!�6U�،"k�DC5�8�8����I�s����^ƀ��-ػ�7V�zfxt�}#S����r�����=���ů�DSz�D.ũB]T���Z|Ư����Q����^R*��ׯ������������(��ӎ�3���\ˠ�r��MK����2�N��Z��>>�c����߆���l��~3 ��p%֩k�o*�s89���&��A
�̆6&E��f�s8���F�J<gvҫ20���;|u�Ə�����k[�$��8[�u��'��:܎���З�Tpq�o)��}'B��u4�8**}�#��b�����u)�����a�bG��u�t��Ѱ���B�7��mS~>�B�+��g���@:��j��f��=���ɋ�'���>_N|b|�Q�f6�V�R���9T������g�8u�f��u�t��o����'O�j�s,��q����jvJ��%���O�{?4M���W�k������n��f�Ƞ��}:�o*�?�b&s�)��0)�/����� �}�o���H,�o�Mi��Gj*(C����u#�|���qGQ��rb��E��:;��۟�'�juY���)��h�������'eN?�gw1L��-LE���E�ZVð�%����A�8K��1����b!%S3��+Q�ݔ ��:�ηmd�7��"l-���ty4���������Js�B��Sx��abj���djQ,��F�Ij���f�$Ks��P��~K��_�`�F��>wI4�����x��|���Xϛ�@�]}Ru%p�e0STTo��pC[�5���׫B+~������eyK�vrC��n��B���L7�m�z�E�[)�WAx~rQ8�b ӿ���}pHb�ѽ����(~���o�#?s�s�_����X4��8�x�A�3SS'(��(`{(��y$D��o�\������]Д�t�#k���+�Le!�}����V=������J52�J�p���"Ou�w�~�S�W�q&'K�(�܂����j
{u:q��+ݪ���?��f�=R�tN�b&%��<;�������쩮䣇�/i�|�٠Y�`,BV�S�\��4/����@�J�o�7&vr`�m_�[Tebϣ�#㊜�����B��Zm(���p�)c���P�L1"����o���4��{�c8��N舀���&��h�4��T��������
]ϳ�{?�H_-50����">��.��&�U�%���� V�.�A1������F��.8 �W�f+�� !�u��j��^�R���eښ1�CB��zDf�}�F�7����}�_#�h����(�?���,��u�W�)���?Û�i��ȁ�%��B����{X�
Y�kʝ����M	�*_�I�g"'C�WWX�
%H5���i�D��PɳP��dfs=[�v#�Q���V Gn�u$�ß�@�I@V߁� �B��t�C�V@�n��xN4�j�}�w��o�;�K� 쌖����L�uqr�^6}�sqX���u�C�8s⿴������Ž���d��N��}�V�v/0��]Q��!fX�8TB��y5	]��ytl]m���L$˳��_���v7}��A1\�MX��Np�SNNƹ]&�>Q�|�@i����L�cZ�qSTY4)�Q4��3|�5��ϛ���}�'����r�l��o��\���ڻ�ϡ�	젳WFS~�\a�Ls�#�q�ab.��DcVAe<�q��-��%I���,Y�z(��m΍<�wC��~v�˃ H���|�a�b��,�����|�D���"��=	g����_1�z�����ag�k�X�cI�q�w�����w���e2Ɵ��CP�.Pܗ���R:�:�] ػ��9g��lh�^���uݞ�����xξ�Yld*��5�$Y���%Q�p�����G����־� �%0Yy����P���_��#��d7��!e�["��<6/�����Q��A���~Z<��V�2,&��d���!�����}E���'���s̢EN���Ƥ���t �D\؈�n�8y���"d���>[�l��2TJ����T�c7����_��=�d���Ol����z\t�g�e�]�R�� F�E�{E����GZ�w�����*�%�qˌ��9�T}����9^������aR6᫠�Px�3|ZW�]¼�d��6���lзtx����[]��2�G��q���w�
���}�8��8M�	�:��Cs(Z�����J���������\�=͟�m��.�$(���|9�Y�8��yv"��$m��H�w�Tn��E~y�~�5w��~cGC�<.[k>�ٻhh��~D�h��'����T���K7�Wj3]~]��9���hr�W�D�kc�=|K#x:��S��N����,�Ԣ)����Z]��T�6�b�XҮz~�S��z�_�z0�P<�"ˍu���t��q�+T��HϾX�77+�ǿ����M�8��s��p���_]�=x����!j_��rr��/�fq�s�"MՋ8��:�A� 1���#��jƼBA.aj>���p�[;?�����B�y��
Yc|o�oWv��JH�	�����p@�*�����?�}p��?F�N��?U	 ģ
���13�w(�7�\�|�{I\}o��s�a��{?��9ϲTW�
:`{�d����b[�f�"�NN�{2���t�'5������;8�^�����iT�8�O����b����;����Yׯ;�9%�Xy�̫�GY�wa�����O�Tg�q������X�t����{�!X3�N����yyעZ^�Q���9H��R�ٍof64�
�&�T�ä�}N�q.���o�t��E�P��j˓a����n��6]:����yN|�f5�z���[u��[*�F�c��"����Otǳ�g�8��gOi݀W|���
�������:�<���&4����X��EV��!c��������R-�V��U����������e���1g.q����N�S;�uRW�nu����E�Tz�R�+�7Xܴ�����'���L�(xE�n��&���3�C/inGJ�A�����(��P�RGGez�~�60^ͭ��Q�[t.ѭ�b����Y�!�8B��r����	h:*���q݅�v��*�*Ǐ�)���j|��Fyu�9𯚼XDt<��ф�+���}�%��񚚍"��Η���;i����a"�i��O���ʹ�w���*��H�1~�ڬ�[Q���,�`l`s��"P<"ݲ�'�Uϲ�����FPβ�d��[���Λ1��Ie��^�O��o���]��/m�Rn� C� �����i��d�&���K��`,!��۝~ߕ���_x�7�D�s��Z�\�>�?��mj6]���贍|���ﺁ�̣�`����^p��{��q��s�IX�c�����!�ѿ#�˵�n��L���m�l�������j�ύ�K��� }���?w�f�(���� U�������F��IՇo;>z�/�jG
��eW�"�(�ē�+Ƿq�1�+,��-��{�v	��Ff��C����a��U�p��P���O3�2V	]���"��F�~Ss��?�x�?����䒛;�6��.L��ݡ1�f�*���*膾���oL}X�28PK�s���0?o�+�`�������d�K��XY������Cz!��8�������A<�nX���@=����*�kab�N=FW���3| Ō}�h�
]Y���>ɸ_?���S������b����V������Y��&x�˼���ۭ��u��ȏ �������Q��Ǭ�a�W��Bg7���s!�3��I�W�c�kc�8�+�Te<h�R�BcU��yd�Rfc}�c�$T�DK�4���l0i��g$�<]ot�G��*�.O}�x~�z5zo9D`�Ġ`�Y�5z���Vt��YԡÄn��Ir�M��1���t�����tZܮ�*���P
�������J�h����Uj���h�!��CL{�:^�C����gl���}��rSr9��N/N�i^HWc�RU�`�8T���龸��
PY���|T.d&7�a��.�΃oIÎ�3 �X4Pm�����>@�o7w�������$����,��.k?��`�Cl��AX�{�3�/l��ؤ��H��0���d-��xy��K����X<B/wް��7+ϧ!�sx/l�Y�L�����P���X'2���'���9�����JI��p�8��˻J��+D�pJ��A��Y=K2p�(��꠬�HX�I�#�[q��l�cܓ0@�?(D��E�П�����A��\Ā絥�����o���8�ź<߾O��c��}'���s�E��~V\�aɮ ��pd��7B���0E�P��O�;e!���'r@|�~����w�yQŏ�N��v4����I*h0>�4�
K?$�ȋ�Ր�eZ{�?$�;��9n2�(vDx�>����䭑f�s��t�`�Q�:Fq(������������d(���������	�cH��W����3)�X8_�7T�ܧ�,AIP� �:���j?a��� ���
`����S��I��"���)(����xe4��|����D$L�n��wn�Y%�����-|�i��\Ďވ�&�P<��`�[d~]{'�گ��1Y�"HY4xm��N�/h%ǁ�o/��.Y�㓲��,��L��Y���3G����Z�Z�2~0Alv��u�9�vlņ����`G8�G���zI6C�b�����{�K�?��Q�[qb��mz+�Ĭ)��?��aq/<�ä���X���I� �{g�h��z��Y�wD���V�w�g@��P})+�l�|a�l����� S��@p����uL�� �������"�뺁 �6��7�jN�K^c뀂W�f�Y��%Zl�2��R��jk��r����<��.I���*�-�Z�@y�d���I(�n{L�|d�8g%�[L����C܁�Ip�/T%Z���NM��2N8�K,�h<�W%��|u���I����â�E��;�/�,.�&�
L���S����t��.���@99q���̡��9�nIgN�Ӷ\�K�'h���kT:)�����#z���������?�g(����et���e[��O+�q����|�.d$�52A7�C�5�z�/�n10�����`���v[2�u�Gm�?W�uu\��E��"�+5��ÜBI�rK��~4���H*�)���J�W)E_نT��
�$�D��$�KF1���������m�))�xq 0~����ĭ���oC���z�* �>��(#i��i��,�~��.���p+��N��#���b2]�OL?�����ʍ�2����G�G_�o��]����mkB������m�%�4"�T[����u}-���YuR������9��
)഍}��[N�2�Mƀ�ˡ��~K�7lN|������7)Rh���Z��d�Ϟ�69cX��'+�)::8���'��y�We��*�������핀�j�Yν@�jYt5����Ǐ{*hG�f��EN:�Sn��ޗOQ}����;��;>1�#O[Ky�hR�G	�]�}T��d��v*�7G�y��z�BC�s�3!f�-�{)�xҏ�tL�@-��Q���bO�}n���.���~u��8������eaw�٧o�Y˾z�2\((����u���Q:*�4�4�y�ʴ�k@�ǲ��`:��q��R,�����I�n��ص������^�1��έ^�bd�
�I�2�~ms��Q�JYN!�Pe�ʋ��A?/>�;tT��S(?���t	5�����9	A�i⎫�(��Z��W�㠒�ā�Y&f��A�`�Ш�LM��P>/�j���qU�m�� �7E=ڭ�>�6C���i��2��=j՜�+�"d��vb�-�B�
i7�=���1�l@s�o>T�y*"e��Sr��!�wjf$%����O��Zu�#ֿu.G�Z�WYC|�|��%��C�����U
&�w���*��&Сe��tn��}�E��	��R:�-ɗ	*�yK���������'� �/Ǜr����L���#R
O�����e�˝��g�r����ٓ�T�W��'˕2����F�B3y#�ux&�M5(6q2��r����*���F�˂̡dn�d��3ˬ�6�� �����I�W�N�����0���M�h���5qr�M�:J�'���瓙�P�)�4{���=l�t1���&���Ԩ�H/�����/�]�,�������a5Gp�@�����j��zꢲf���G���� H�|H���ӛ�	�~2��5�ɺb�wn)��(��
#�륈�S.�6�>^��n���(u������kt+}��M���,>
����,(�{9��7�K�YW>����ײ�Z���):�)�W��q�5�L{�`Gw|F�X�E�<��yY���=�L"1����aR�m����a2J'�����Su�f�/a�=�c�-�q���{�� +7�_��.B5�7W��@]���G��ǡ@�O �ON�Ĥ����'����I�����9�V����C�Q�-�-� �������0�v
�Sֻ�q�����˪����J	��c�f�!�J�-N��`����v��I������&�1�'���
�M���{�{��]�o{Ȑ2� 
��N��E�Y��t$��x�N��<�A����M���/�ػ�L��>�ɑ!J�n:�--e�rm�3�O����C��y=H ���jdR�ϻM�9_���KMf�k��i���I3�V�p���r��p��D�ߡX�\Q4���kOYY�r࿝�bZ��F�lU�i�8����9;��.BU��[�$ w�42W�٪�&�+�s�J��#�X�������f�/��* �UC����Z,U�5>�1�w�n0^�O����[:*=M�5\h"m��J�e��++%��t���t1џ��d�\S�ȅ�
4�ԛ�`5Nb�G��LP5bw�������{	Ǜ Y�+���q��W>�ш�Ox��t���\�d&�.�ۦF�iab�dy.$��B&m#�*��q�b���3�2 Ќ��G7��AObȝ#(-X�3��hGt�UU=�n�r�ƀ�����_ޠ�ℨV>���v�ة�[J��)� �-�_˰7�q���F���L�2�r8��jd����3S#���	6�J)тC���?~����2���ڱ���W�ŕ�ߟ- �M�vQ�-�$�k"���dc���V�ˍP�q\7���a4g���ptk�8_KX��6_[�8e(1�/,ԙs�p�BB'�_��g��ǡ� ��c-��f	E�A�� �@q�t�&��6*f���vq�鏌�����lن���У3����{�A���
,�aG7�:�2�/|������Z��ZR9��C͋�����êO8�X�K<A���Fp������,�����5P��V+'���(O&�bNhP�d�6�@�o� �y6o�-��iD��"��{�-E��\r ���ع�FHe���O>|�טG2���s�D>_�u\�_��A�,^��n��ĵ!ff=���b����;ۮ� ��ۯ���P��Cž�WӮ�Jt�	�R[��e2�]�_����h�WU��6+B6}�<S):�m���J�2�?�>��A�ؙMp巣��D�)f��������&I�ר5}�h}Xnu����G��ߣ@.�(7x	�4���'��p�:t�_��q݀�4D�`ڕ�(����RW;d�̌�yX���hX�ZUP4����S��)ftY�4W�Q:��ר��z��"O٢��foo�����y̤c��
CW. �����!_
�+��j&����MΠo!ؖ%��Í;xE;�&3�>�Q�e�II���>Wi�Y\Q?��μcukS��es�wS���z-6��A�g/9�d��N8zd�~hٽ�xx��@���@�(�/��P* ���\���QWWd�(D���jХo���ػ��ms;�����A�����/�98t/�b3��Sy��E��jo� 05�AJ��l~���okuH������p*o�سﲜCc�1˹����ǿ#W3Ks	�"׳0ww�j9���&r�B���hݚ�D����Ԓ��C��"i{m���ˈsYlW��d�N4_�9��KqX,�x�49"B5����N_ʹE}�c�b� ~�#K��C�RU��w��
W!�x��p%=�9B<�a~��r�v0Z��29ۀ��ER����F����
�؃��4,���ߺ����kKx �ŧ�$H-@0ݎ��܈����=�����nFO�A���d���7\?j��y�
��8�̆��`�H��������M�@���m 0jd�@��	���� �����ueE|���ĝ@��!*C�H���'C���q�a󱽃l�V ��he�j�E��Y�*Gc)�.#�?X�O ����"J�R#�߶(�K���FT�/҉pOS�t#)K�T�����l�I'�WY7D��x�iC��M���>]!���P���z�1g��4y��!u2::࿍��<ko���`��l4��
I��d1�0Y�c�S��(�\�J���W@�@
3� ��'��^�k�PßX���X( 74����f��N'�ۍ5����L����:\LN�j��X�rYQ1>�^MJ��~�F/�֏P�L��kj��C2C��EA��m^5��q~���!����a����Z���ӕ��斥<SD-�f?�r�nZ�7��94]�B\:�2R��,k >3�!$T���@KX��3,���R��p�����0�m�:��fK��c�Y�����B��0�^��x#�!�!V�_��M7�|eQ}n�w;|5���kr�\�|�x��JAE�C�k	�C�:9d��Ԟ����I��x0�B �,���vÆ�sX?�Y�Y�v���O�f]����:=/l�x��:������;��V8E�S]�j6�W���y�̈�F,O���+�J���B��F����C������p�E�B]��$⢎K-�Bw�*j���I�YUJxK�����K�x�5����;���|�ߤ�M���ݜm?I��l��KԝCp�X��l���L�*@�����e�楎*�l���QPsl���_��;G2�'6C!�w�|i��շ�x؃��%6o~��MS|��m;�J(�D�H�!���B�m���W+�\�Tf��Amw��K�2��|�������"e�,VB���i=T�G�%�J	4b$���2���@�u�)�_�4��9t$�x��K�C�ZJ��+b��?w�pb����wI<-�*�	Ke�#;�U�]֡��	(0?2�a�i;W<j:�X���b�+�t���e(���i�GC`>�m�$z��<V�su���ܬ|�w�L �/|�>�6�&h�8:Ė��qP΃������1*���(�0cx��K$%���%s�N,��xHR0K���z��X@c%��O��LB:�%���(����f�>����Dbe-S��(y�?TN��!?� H��_��r�}$�Lg��B7��A�-�F�uW
���Ǩq�@;
̶�� G��j���W�&4s)r!�SiL��	a�M�U�k6C!�9�9�O�/#�ҫ1�Rś�{b_t����y�ʡ����C {�;?YTZ��Kc��!�	�/&�5�x��+���6�k' ��{���*B�Cr�ρw ����:C@4O����iI���yȎ�Js�"�c#�Ɏ��
��r˻����2�����M��_}�j�cP,�/�M�J�IH+�G\�\՗С�YF�R8_V@t���uE�O��eD<6��'x]+�d��,�&Yp�x+P�fN�̡��}�{�{����&$��,>�����ǋ(.C=J��|y�c�y�?�(��eu� W���4͑��	�<	9�����1i.����������_7t����uYZ�׋thG�}�&ȝ� i�RO�y,ܜ�����~��E��y�F�/,���K\�.�������Lڀ��A?VJ�W,P��ሴ���� Pk�T��uH�(&`���2h�cCH����w���(��N$�	F�������H"�n����2k�|=��u��j	�����fT^r����w_����%`�������P�WL�@m9f1��ͪ�G���m�u+��EE7�,�T0O�]�Z�v�`���i�~�|C )0b��!��0|�" �o�ʡN�R�,��aM�p:\�O�������p��\���$��q���1:�m3=_C��Vg�����  /9�'z=� �	�=_@
�0 $�]_�,*�6��eQX�K�^I��������dYol�:]�9��������8D��,~�G���3��S�ϊZ��q@|�0Q� ���}t���Q�����/m���r�uv%B�ri�>nB��� D�ģ�6ߢ�@N�o�s�f��MK]ث�#?��7*ʱ��y<���I�0��0��·�;�㆐�|� �����,��^@UC3U��4gn��K`�*��Y( ������y��x#1HtAUbAԔ�&�q�{m�8(<�{sH���5����a�ׯG	�D�e IUy�<�NP�q_�^���zZ
j��/�UV�[�٘L^,�윓)���3S�8>�Q���T|�0tEw�V>*nj
���iL�N}�2�ɿI�gL�����E4��	ȩ%,~�3(Z�bR��/��B;���X����\
c�͍�#��H/��?&��B���;�4.ĺא�`�,�s�!h���@���W�o����׾�c��Bѧ��F��C��Ƌ���ۼ�$K+uAo�}��įtA�#6;<!?������	���o�!���$�t�B�)w�'6��z��ɏ��R2`�UM�b,A0%�@������nҋ��>��Ht�r�NwԀh06q�:�r"�Y���)P��Yqk�\1����>��=�X����.D�����\v _��кɑݻ�]��
+�#.�pǛ�51S�u�S娴P"9%1��m����P'��&i� vv�Y�`C�R$ 'W.l,C���w,��hu�g�>��4RgpS��bu=�"�
�8[X��c�x+��ڸ��*Ǥ%fl�vK�* ��r_߉E�c�2����=��h���
��kni�'Y�'6�|/�&\x�����+��];i��}�|M䷧�aȑ�t�n\�=3��CX�.��� up��(<��:�@g���IigjP�ͳ�������ʟ`, ��	ts���8&��w.����K�a	ͬ����g��YGG�O$�p68����r��k���C�*=59��;��sL�c_c��e	��x8?/�����:[@��^�a�$ht��HS�cN�o�����#6�&�h'�\���?F�c#7a���}���n �{C��+���^�(�r�X ���h콻!��!���B6v󓞟��<svAy.���-Klդ���!��β�����O���p�{6{D>͗Υm��3�|���YAq��Ȣ�P�uD��i�Ħ^B�A��\��- �)�|�'Zl���uL����@���p�t8B�/n#�b��x�(M��r�YOd[��KS#��1���۳�i��ށ�-r,$%hw��Ԥ7!����F��Ua��G��~��S����!kEK-��!��B�-! ͆�X��RM�گT��l�; �h�`��ի��k�n��K�榧q�v*�ʰ��)S��W�W¥,�����ީ�|aw� q�sٰ��t� R<�e�V���yy�s��|P���5{
H?�����%V*�1-�U�JJi[��*M到�x��c�Θ�ʕ������|�x�'�S��o	�7���YM��s����kf��j� �H�]l�3��C��+�1�����j����������G-��}	L]��!���J�2��/"�6�KE|1W��ũ�G��"�-����%�3$V�G�.���-y��D	�y���CѦ7���xd4k �ۈ7t��w��
��+�G��(G-fi�/�f���@���H��G
� R2��h5��9 ��6P7P��Ѐo����m'~���W$$)�u��
�D�0vU�ý�9�yj�g�r�wO� )Eac�?�>�Xߑ��shf���
�K��J�u� �pM~f���j�'ɫB=rX�4�s"��u�|K�e�����k�S}�F$�+�����aE'f%e��y�'�S����4^<�\����t�|=��p�G�=q�"=���S�?զr"�E�IC�dq����9@�M�mUkO�ԹM뺕�B{���H�:�L��n�Ef���e�����_�5)	�F�d�?��C�gD,]��Ƕ6�tVw���[���6��������H�$�oX�r�qI`���ç.e�Ʋ挍-�w_9���;�^M�Lifa�/�i�#nRH�-����ѓ��A�[���J�^kC$�]�
=�7YWLUӘ�a��oe�b�\KE�h�l
��jV7��(gV~"n��Rn��W�H�ֶE
چ_2+)���Ij/��K���t���Y�\����Sg=���|�.���+�է.ٚZ�7k�0A/� -4�i�mV2,":_�������Ɗ��kf|�*qw1�y�:�r,��v��ݔ\��}�P����g)Hj�8y�6^�e�-f�9:��P�vR:����@����hQ �_ډ���4�Ц���Aj&ס?E�e�j"U�;џ����e^�`2��8�*b�Z˱�$V
���K[�C���!��>�ޤ �+7ܿ�Y!=�P1�:��{c`���ݭ�]}��[B5��H�v��ԇ�t_�D��@�lQJn��ŭ
��R�Z�����W�H���-���OVU�֡����BPU`d�|z����8(���0p!/��ͫ%��a�T��af�Ӹ���aW�����x
���ul	��l��&��z�7ӏ��*����k��%!Dk��|��b�v<o5��M���e%���}��|�&Q���>6��ئ���@zM���\�x�ݞ�9��(��,�ߦ��]e� wц^�D?o��c�v�Ґ��h�k"P/�7�v����������X��)�D��7��tm����U�˩�|Ǒg£�%V��T�}LT�xB Am��G�-�s�
t�:a!�$��N�Q5����c�$�c�a��'�3vx�_���͹e_�B&a���>�<߶ P;52+iL�ׅ�N�:�;�J�������%;��������ZNn�c=���3���i(�� ����� �E�{ns�K׿�Y(g=��3�|�X��;tK�ǡǪ��<ou1��ܟO"���][������l���G*X|��pZl����]���z��Xq�N�ٗ��%U�?ۨ��W(��ܨK�k�`~3��6�czI�f�?5�^�튮:�4�v��9`�h������{����C�d�g��+-�yB�\�N�`D-.�>�Q���D����TKKc�� d��H�Q��n��3�Tc��R�r��}���u��h��ݗ$�P���V���?�ڝ��w��ɭ�Y\��h����V}���������P��"�
<;pq�4�<�#s�G�~�U;xMqҁ����]޵X'��{�*�����5�f<&��ӳ�.�{D�ߕ-?��@�9���n�$<�<�4!(I$؄��XSS���<�	R��R��B����rX{×���9H��츊	�������{/��Gh�@M�T�cN�X|�@aߴ�����	��Z�{��L�?�0�O9�+{ɟ�Oph�)p	���h_�bj���2ϜȠyab���c�)S�L����+�SK��V�Ч����;������)��%�z���#��5_D�l{TWk�g�G�罉������e�.u�i)qKQ=h��3�.F�@c�Y�[t�O~J�R=���4\�=�~z�J�x���� �Ϊ!����֔�e+3o�˃�`��͍Q:��\�9�^��2 ҂j�vZ,h�(S�� :La**�>0�8�#�D�nn7SD���Ֆhq? ��,�&��,�����?A�W��,��K�i���km��n(�)�L��ğo�68�KP?��+�Lݨ#t�*�yv�d�3��d�oʫ��5�]���V|���(gbJ�!b����?�d�$��b�.�^�$�;��Moj���C���퓝 �pLr�r��%�3�6�L��� \��,�n5��h����]���>6�d#��%�>�3��+��W�;��O|j�R}�4��[.8�bO(rӺj����S[N��t��O�M*rs�ʖ'"��Y��[���%WSD(��uocqg�L��THP��ia$3���ֱ݃BI�n��H!^�㮓$HI����iP�$��sBx��{1����{ϛ������}��gR���k���7����ti����N�X�� v����3��@��������E$��e����Ԇ#zY��=
�8܏d���[
�?�D��mY&��dD��4��ob�ί����rHx��aC~ӯ|Sw�eq1�~Yg>��uMy��׾�,��lI/�6f�G���I�Gdw�����z^����w��mM�r��T74���u>�}�o��	���X����Z�9�SǪq���V  � �cj���;dqݕ�g����q�hA�K�`�\����i �Q�V�;�������04d�X]/��I9�x�ZK�w�	����&��@�k��$�>8���P���;�{��b���8����0��+B�.�`�<_�I��}�{�9O���7Y³�/�8A��u��)�p����2[�|ۛ�A�Vɒ)z�SL�<�;�� N�G(1rp`��8����Z_�jw��*Y4i'���Y3j:��/��$�-�#*�� ��M#��޿0��7��[����)��W)O�h2�|n~0�|��Q������R�^r1�~79�,g��O	�ykVL'��c�ύ%#A�	z0vF�Iix�392�κ��W�;M�d9���4fHX�x����Ɲ���L��9�q���F���v$CSO�+�����;3K�6X^O�v�ӷ���E�b��א��8�աc�OOlVϭI�,�	'C�5��߇J��2(���e�͞��:_�r��l؇�I�Qg��,�3 ]J=���
��UƏ<��xټ�f�IJ����R�d7��9ږ���h{��δ$�SdK��<�*�"�S"�A\�e򛂖/�3^ h��+:�6��#u�㾱�y��m#��V��Ұs��?mlsv �t>sQ�՚F�ޗX�/7�;�P�<>�w�	��e�&��H%{/������(��B�__X:��ಌ��0��xȕ$�cI����bJ�z����Ç3�k ?}�[�@΢P���fe�?�*�@���R�Gw�.e��RE@�(��f��9�S̻W1���}y�Y
Q�xp�:���:ڌ�_�m�'��_^�i����Ѫ!��n�[6��?�
��H�j4��5�?�� |����7,}�ʡ�ћ���E�or?<2�����SQ�=$	���.�cT{�{�~�X@Z��Q�)���E�-dO���X%��x�W��<���n0p�$7�c(?��c�����}`�M�_^���Y{ �ɲ�V����֔��V�c�[����%�]cM���7��U\^&rZ�><��X�$��V6~�k�m�{���I:L@f������V���	JC[[x��B9��7-�q)+����g��;�PƊ� l{3��^�yo���m�!��8�Ɵ|v<�4 ĭ(���*Wߑ�dnT��Lf���5��++.�����oR��:�þʢn���0l��[���͏�/V���w���6gx�m�	&��y�[����k���>�g��a�������D�1Ϊ�0�?�j��n�Qf�w3�ʮ��!2%Xէ$��2 N�$X,�����[G܍�W粆��#��o��J�ܶ��Fv�R6UE%�3��<����0e����m�y�U�Y���P���@�{�!{�z:N�@F�9g�H=����;�]���(<�����N�Ge4bQ�I�����5�/�H�ۘ��A��Q�h��@+�T��v��wE��f�5��-S(�`��r0����8�$J�%��!�*���S\M�5:�{pww�w��\�݂$�;�݃Kp�!��������?�V�S�JR3�{�����9ӃG=|� ��q� :�NǛ����Fc0�f��>$9#J_䪼� ����9�jғo�M[H[�L���>ETs��Q�~> l,-���/d` ����"�oкՂ�,4���#�>9~� �Ȩ��mк�6�ҶF{[��K[�/��G���ɭ��&+�N�E��yL#F��r���R݉'4��&�j���}iz���sił���3�G�. vѯ�?!�����Bf���Z��{W�����z���:Y�t���p7A����z�1�8�&ǩ��t{c
�U��g
���.16�0��Ve�����4wH ��#O~��u���F�k��ل?����p�g���1�՜�_$!_�?`���6���[-x��d�z�ST(��%^U�9�&�Lw��Q��1�����&�:*=����������WO��exPv�l��ޗ�CT���xs�op7򴞝�U����M�x�~�z1�����JXFދb�'����Z$�t�=�`]�}RwG/�;��>o-���)ԠyY{�]�LY���ވ�R=\�0ZKV�{mkί�o'�c$6"|YJG�V��[��Nb�L��B�sV�����˿5[7�E_�G�`B؟io�(���~n�;Ǥ� Y�'���~�Wѩ��֒u�R�|��i띔�D(h��C3��/O"D�A��ƀ�5�Q�PzS)�`��	�<��\!�K�p���^�m� �Sv��ń�^g�N:#F
�jy��;W�%�q���X8�&#G�@x�F֖ݟ�O�Xx�V~Ub$�h�z-I"�$?{}�x4qLˎY�IC���̪A�h��<���ѝ���	��q������i��2`B�h�1&ˎ�笖?u�*�E��!*�Bd���J�W%��ʬ���=����lR_��ڴd)��~{��!��u} ����S�ma7Tj�́<�F��d��l���IOJ̄����;�6�:��Q��,��S��Uo��<�6�~�	L�{J������UI�g˷�qId��_п�¼'��`)�����!�u�K5V<i�����m�!n�������J�ۛ:�(�.=_�G*8��E����rj<Z�5���6xr��iNѠt�SҪ�����&��~֪���{�F�P���Ni�Ռ�^�G���Y�ӪD��r�z!� ����D$8I��Q��mKY�N�-�B��ā�V��\$�<9�̫_��C-T�5�'�BYao�޻�͸}^��x�{Pw}�*}�t�T���N�L���Z�����E���*m�7�����ᤵN�)w&����{�}��;fU����6�%\��9\6�Dt���b����j-�.:�2�V��P�F������<g����)�A�!\����ϔN�\���`ժ뢥���4:�9��G����/JbD�cbH�&P��W���D	Ŗ���JJ�\�F�F�I��-Z����J��I�k f;�Mo��>!y�`���TLf�>'�94h�lP������E;��gT�"yf���J�z�/����)�N�du�7�����;�YFX~��R�҈���4&��nq��T!3smv&zf�����:ܾ>�lJ��JEc���<s\���<'�����H���xc�
s
�Tm��$X�0D��;���&�Vs��?��$%�lV:a&����>sb=��=z�D#�Yj:�d+�S�o�~���3��;�,C�"b
�]|x��e蒗���%�� EƂY���	>Y���a�e�Ņd�6����7�g�^#_�����t��m��[M�Q=���A��	zOe���4�V_T���3{�i��4wC��Z�"э@`_
�Y0�tur��?Y�<Y�֖g�L����zy9I$��/��F�9�����d����%lxNo�=����W�T�M�ǎ���h�1��@ҨR_��f	�61����y���=-�?�&��rV�h��*�K�:�,�^?|M2�mM�� �V9v��ѫ�*`Dr�������yz��Y.�Y�W��x�&��9�w�0K�ռ2\w�nH4q�Y��
$'����(Z�V�"QG��2Z�5Ԕ��O4Hw�x^��LZ��I\JRz$VR��:�����&���������]�����qfT�(��$H�Uڤ!rн7�A�X�Q�۷+�����Rj�đ��>��H~Z��e�`��<`X 9%�~��? ɾg*���S��H�*w]J�ND���I����'�m�)��A9ip��JL�h�Ĉ�����%>�y@@:�4/���r3@	���\+D�-�D[y��溉;���Ut�9Żp0ɵ��R�A�S��ʠY�����]k�ߍ���w��.�,Wä��g�ǚ{~=����Tۃ���h՜�>L1��.��B�l`$��5D~L��F �w��)]z�3/Q�����\��*
$2�n�*q5(�4S���|�2�Q���SX<���
@g�OU_������9�����G1o�wp�u�&iC}�ar�b���L�wT�1�Ñ���t��ް��c%O�~)���x�>����s�F%�*�uĹ�	��(���=��}I�MFy��Jͬ�A*�,W?�����-]��$��'�$�l���k �e]J�1�rVl��w ���a&f���ǃQ��d+Wĉ[�V�ɽ��:j_�������}���x�"���ϒa��F�48�Л�"Lv�6ō(!��������}-<��,�×������3&l
�j����OY��0��o枾�iYSY���hm����uѦ��G|�1�+�1�A��y���Gg.���,��N��=c�S4PP�1�3I�����ͥ蒡�]�r;� ��z̲�4�uF{�~Z*܀b�np�"P<'���'��R����e��	P��O8������W˃N뜺����ä���Q���_��m�7�#�lf|�&v	I�%����Z����)��N�!��sn�D�rS����Z,��"��:?�`j bh�k}RL��>��b�&������mj��sy���9�z,�"+�7���12,�K��-@�ϤM��Ҭ�
�bx�%�W� ��P.��4��=�؏��@I���Ь�x(-��眄[6��F2+����Q8����YaAlC�\�L\"�=/�w9���Ttdz�ɉN� ���Ҥ��4.{1J���'w=_���5E���Nw<!��f����G�k�j!���2ǒ
�Ӹ4Z�_(�]N��
 G��+QN���y�X�O�!�\�2V#5N&_�іo�0 |�NEl��Y��4�$��!�*��
�b	3�����P��G�v��_�!��͵tA���/�/�y���k^��:
%�T�J��.�h�z��Xڄ�#\�U�7�i�ʵ����J ��m@���U�e	���n�I��;���z�}*��s$�º�La)��� ���|ǩ�#@z:x��}�ϸcZ��LB�Z��iZ��2D̉�^L
hOd���b$�
����HU#����d�tW�.�4���ezسY���I:����S���ضke�(��a/���1oj�]XV��g-K�_ِ|���D*�Ts� G��f���Ӭ����_��'�֫#O�za���.�h�|)�0Qr�g�K��Yx�E�ӖVd;Y�s`�aRhA����AZ�c;ЮV�#eD�o�J�+�|zʨ��Ө����*�3*N����L��=���Բf�aY��نɋ����Z趣,�ɥ��OMȁZd��m���c����tBׯ�F��p����Y�q���z�(wV�O^���+���Xޣ0˖=��z��g���6>J֮`9��E�qU  M�E
?�I�2��yO�T���m���(� ��r`gk)�Y�H�j���ȳlB��^`q�y_��ih�-WCa�A�	�z�qav�*���qj��v�DS��Ng�h$�� F_��^��6���r1tvtY�	P�3�	�z8�{�
�ś�c�q���ì�(�\�=T\A��t��O�L��?�d���?R[�3@Ub��)��R<�S0�(����%�g���Y���IC*i�lד�Z�V�Q����5I͌U>}��9/4�#�l�c]jl�{��%34�P^�E��u�����cY�V���a%�ƃ?��8��'�RF�;Яi�^/º�m�zg]�Ty.h�sb#�J�Ԝ�w��d5�>��uka�O�I\�崂���ia�4]kζ�'t�%��A�r=���(mX�	�ș�o�0��7&��(սb[�� 8���0Å�o���|2��8w��=��)kD��I�ŋ�d�����I#+��ݽ��e�����k	�͏�@ar6U�a��x�ìv����iC�� _.;�9(n��Y�ʧp]��Οk�����6kPh�"���V���:/Z��i�km�G!P3XX�C+�{�Ї`ghh~�d9�
a��%�q���?NR%W���1;8���%��A�����W��������x�e�@�C(��k�a�+��+����d|F�f�LO����Pg7}���-��èF/�FF�_Ү����nis�9QY�f��M|��� ���Za��G{����4����y&C�kmM��4�gF�iZ̮�k�V�Ƌ��7��X�4�������	J#¿C�������1����:�Y�<��P�7��O9���׺I�9(C�0���vF��
��$�}�8y.�����3?3��٠,�ph�Y=-IrԳ�5Z2\�#���6����>�����{��#Ɏ_ln�@�R����h3�?���_��[l}�X$9�������o��=מJ(˔7^2�>m��/��ԿV"I|gv~/@z�? ��ME�b���h�"t��P<���`y����ꃊ�w���e��R.���ŷdmkd��  �&���.�	'
2�b���L�{ꌧ�Y���L�7�(�ZpX��%����p�������f!����a�����O�/�����8�h�ߘ�Ja�|�ʗʷ��s�t�f�܅j^X�)y������NHr�<h2�!�w�+b(LDG�%�{Y͔[��~�p�\�2_�:%�E��r�S��lQ7*zC�B�����&�^��G����q����0�Fz��7�F)w��0l�GY`���z�R�@_�M�0�S;�����5Kȣ:�òtK��;�h<0�Y�S,�U ��(�x��P�&W����>r�mVE�ᨖe��f�;_���Y�.1�����R1A���l���G���|�as���[���h|�(�ը��܇�\׎��s�sB�9�]�\bS�l0pWf{�}��"� dF{�G�]\���~�N��#c�����Q���e��*��z��w���D5uE��f]=�W���6�9Y{�jo@C�8����������)з�:jg΀U�;��٫�î�
���ӈ=F����$.� �Eq��[�������ˬ=��0<��O�&��-�׳��7��w�z<XI�������:�@�Cݠ\KO����:���b�g����QO��c�8=@1�Š�.�H�[["ӧ\�����Xq]\&��w��Zw��7U&�����^0�xK0�'<�c�g��0*T��,�9��ݛ�P�4Σ��"玺���(�"�'�f/0Ѽ��M�B��p4��<���iR�����
�a���ﰝ$%�Q��.4���*�3�H��/?�ԄI���5�y
<��!�֕�;F�4���D�,A��FK'B'��S-�������>�ǁ��韗�T+����t)=V�S(G]	ͮ��+���4p��֐nB�X������n}ģ�5�J�Y���$E�������}�4����D�t�Mo̪5.��o�	l+/m4�)�����*�o����Y��P�'��$dJ�M��	�e�jN�x9ܝ=�|�QB��zQa�˂LL������c1��O�����`H�-|Ș:���p5�������}(���V��<o���D��@�n�|l�ykRв�bz��[
��'ʹi�=I^I��HV��J�ne�9y'r4�ލT�D�D�h���a<p�[Zz��Me��Q����]��{�O:��NφEX��ʺ��Yǂ����Ig���N�T�'��?V��������=��0A�;I��!U�{���/�^�d���2��r��	[���<���G�U@�i�A_;s�EyrVh��k^K��x`�?����:JF�:P~m8��`0��u��d�/8�a�ۨS�&@㫞���F����7��r��d�^�bҴ�!�,�3V�	!�w�
U�B!SL9��p��`��a�����i|��]���v�ߛ�P7�%�B���d�ϐ���s�A�8�c=�Y��ň�]:ģ3/�&o��0,�|�5�_�x��1h���<��+j�؅͠�,o�-��B���cC2N�B,���%�)ȅ��p�����FOv�s�:G.���I\�phYH�f2v�0��D�W�l�V��Mq�`؏ߍ$�n�/�W��>i���	�ϫ���R�?z��؜�[/�gx��ġ�v*�:ѐ�Y�k!t��B����u���l˖�h�s�5b�F�J��*ҟ�i��g|��c��ײ��Z��h~�<�<�;�����1�[�m4T83�""�h�i�'�#�{GW;�����G:�+mZ V��T�����׻]3	��ĺTZ�N�2�d"F&T�S���1��� ���r���=c��xQ��d|��i�z��hGt��Hd���V�M���l�հ���������K��C�.c�C�T��0��Yy�6R.��$����&��Bs�D�Z_��"��ڐ��)3;廉o,PS���T =�	 'L�.�k�Ǧ��:��\t�v�V�Hg/G.��ځ�&/�h��� ����J����`xQ9�F++<�xc�{��懎{�ጓ�!���=��u�ߋ�����,�Gl���CM���L�m�5G���q�m����`�Ţ6�He1A�I�6U��@p �j��/��MV���G�c����N�1�h����)%��9�no�coR]���@�xR���\��j��}޳��rW#e8����z�W=o�6�Y'�����[`N��P�x~xI�����Y]-G:O�~u�_Lm�o�Xќ�b��������	���
����P2���������\3�<#S�Jj��d�EyC{ĊwW��'K���e������(��?���V ��/]]u��v��ygy]�'���O*����q;#Qv���'���]����d�v(���g f�>��"�[�ל��!��d�l1��d[e�&�OQ�
�g[Ggm��T�(����̹~��;��cf�GO���-8��a���w��(6����_,����R�<�P�a�<��d��Qn�=�@&3�G5+}�2�B�n��Fط� @凮\\��U��!1b	8CUd��Oa�|.<<8A��o���q�(��\�:\^��>$���|]��N��qSqq��#s}�PP�x.+�b|�~3G����KA��+Z�G/w6��B�CR���&��d�}O$�Ǧ�i(�z�@��F�V�b)�'�i�C��*�������F�j"�:�!(!f@a\�1��O�) t54R�B��B��,{nB�u���3�/�t�2�gǐچ����z�@�:��=<|�k��{�SL*C��uz�l<��d��ly���y.�Oٽ�&�GL�gm��@f��p�Z�b��&a�؉K!��JʕB�\!8|MTG��-w��w�(�`rm҂�_wk���A1hb_�WP�����'��3��O�GMt����>�@����;��*f~d�g�j���P�-�Xҩ}s�M-&��@����$̠��4L�Z>����G���[������H#2f���f/܃�r)��THuH����H��<�:pzT��[���XVRd�NIm�6�Y<E5+����s�U��f���Ay';���l��H)
&����\p%��L6o��F֩����m~sd�Ќ��F��fy�ͩ�p�����͝Hڻ�޻���m��o��p��p�t� #_�?�U����������<��PU%4�>�����R��^��Q��;���[���X>�3¿R�oV��z��F/,lV6�?�Q�S��J>[_���#�N�(����nJIn��K8��	c��b���ħƉ������/$a��/M#zOҨry+�w�a�4pf��~�7��9!)��8n����S����l�8Ӷ�n6� �\:!-mA��v�T(8��4i9�dBB��QGb�b���e�.�w��kq2�}#B�b��׊�Ȓj����q�&�GB�o�e$�Y�������S[P<�Sš��9�J�����u9�n�⦾�(����<�
e�����gb-2��l'�P�5'�p|�Nڷ���]�c+���wm��
�M�1�u�;�v#�U�ț��%���.\JԦy�݇����5�%#dy�e��F����a/���>�cnǂ���>�q*��
B�,	}3���ϱ�1M9GSegɡPH�[�U�\ew:*}�Ж��� jM~��+�ά���
���P��p�Y��&�"E@>���f���1(�Y>��6Ծ���{�>���)�e�ba]��@��D�����%J�DJ�]Ҩ�����>��4�h�M 
�dL��b�.�����Z wH����;��.٫���5�|J��J�;z�c�d�l6�7g_e��0R*�3B�+(�*Q�"��Ai"s�Z�)�g��C��S��Ak�R�x��x��l�!�U"=���w�5{�����֎%��5�V�(8� ���;�=8�6l#I�f�	�s���B�|>�2. �͍�C/3i��P֒�˹�QiX������zO�cq-�++滘�~��D�)�T�`�J�������%�C� ���,�P�9�l[I�!ې���7p���)�Ȍ�&����`8���Z����n~�� [�_�
�Em��Q��<U)��Q�R��Qr"QZ��h"�Gj��.��
��0=T���h�yB�KTow���~<�QŻ���*�ʋw,�����$�;$�]^J�P�|�s�πds�X��1��>e�(����n��h0���B&�F���煄�z�'zv�k(?H;����w܆+4B��2��	�}W9��6����5�6�8�/-�9%T(%4��B��e�����N�C�^����s�	��$�r�7���R�^CL���.t�8�-�-�\S1&U��ʑ���%��3��M�`���Y]Ht�& RtS?���4�ݽ~��ZO��\c� }�eC+��\~1GŻ� ]�a\�+:9k�v��\(�`���4��֒�d�,bZ�6t�bdK��w�	I�tFW�$=���=15�0X��]/�;�eQB���V���~.:%��k�[F;�Ѥ8�5]���߸�.lt�����t�q"%�CD�CN�>�n�t��晕�`v����������e��ZFq�qpao�j@���?P�%@�S&��Âz3��d���3�ϖ�9�0Z��+\hX�(P����[�h�!��E����6�e�;n�����r��e�� 1�Op%CO�2yT���V{J8�����v�oѮ"�Rb�V�s��_�u��R�"ǋp�C�NST��Ȃ>�n�U顋,9F�%�˨[J��_�_����w� ��ø�~��!��b�����Bh�Z��|<A�@��s���b�~8,_3=Sf,���"�N�f�S����9f�-i�w��8FS.�_�xx��ۆ�.4�	f��6Au���n\%�=��;,TW��EG�L`Iɜ#)�ՂY�����.bȈ�����X����3���`s��ȩ�H�%�����ٳ5I�j_ś�]XkQ�0(+��9FaCN�T�����rm2�
ra9$[�ѺϏ�s���q�z0~N���X��&��a���SʿxBrܴo_N9 �n�	�d��J��o4,�,�17c� ��a ��� �w�D��M�;Ƣ�b��Śk鱯/s�8$_v�`���W?� �%"�/���`8�~+~
���ڤ�Ʋ�/�'"��y3�<����r8�'.�^���k��b���ˢ�~j`��"�K����F-���Y��9DB|>m�d��|#,��sG���<�?+0���)���@V�+�.��
xKV�r����ixmt,����B)���=��/]�itM>/�ɐG�$�7��7(^^}[��{�id�.wPU+�dY���]�i$��/�2r��>A�ӐA(���*��m��tòBN=����	���_�?�E���tDS��.�u=�Z@�/�ѥ�?�g!]l�-/�� ����atx�������?RQ�ߦ�<����A��;�C6�tB@���H�[��~�,D�X�4���_82���s��r-T���*T$_OI�{u^n1_$qw+y��0Ch�O��1��Y�օH�|i(��mA6�]���mif�_���N���f�RY���f���~0{.��;0��c��{c-��
��\k4����2�j�(� ��9>p�p��G4��D[6���0��K#��D�yu���?u@��J�i��V�d�n:v,�;ϫ�������@iL \���(}���Ŕ��;φ��I�s�m⠙jfw->.>����>ϫ���٢��}�>>|�	�- �P��k�4������E�� BIӝ��pZƋ=;���2=$�{��� �ẉi��M�.��Y)9��EZf#�%P�����$Q=�bc͞���\E��G3����e�^��\�c�sF� �ܲW���T@�sK~�~^�e� 4����}���n��݈o81`+� V�_�|Iu2 �ZΈ�ͭ"yI������V"��p'��	�0{��s���].�3�j⋞��y�u~��d�?��&1�		��V���+�j��m+}a��h@P��EV�7Oi��k����村S�-L�5#:��� G�E�2�FY�fl"&���W��V$zG�����u>X�gß+���dd��-q ������ͣ��p���Ķ圜 G���'��c�R�Ԇ\�"܌z�VtLk5�iV���{چTr{���Jg��B�J��o�'�ͺ*�����g���r(��`d�kvV���B
���<��,��ZYRO ��H�ʰ�����|R��}�-[G*b�{J�p"��:tw�
���Au`�L�wз恩z:Ծ�
���'�g�X6f�<�*�q���h>=�]�;��c�弳ʩ����4������`�����W�V���m L�V�sB���p�;ܦw��5�w�mWx٘e�Mߝ��4�H+�~�l�I0���?fC�ܴ�F�S]'��#��ί�gy��D��ߨ�q�g�����Ε���$N	}� �f��X���2p駫�_��Pj���ըO�cI]�����cjm�_���(n���C��'���AǱ��=x�����S�1��k�n��u�5
�k��d��i��ýNJ�,{?�����z�8ıT� �x�!�@���X*��	�lgƏ�9�n���@2X@T&�p+2b�Z��E��E��g�+8�}#�Ȩ@g�l�{̸�<A�����ʹuf
s�t���C�-S��]�W���!`�;���@\�#2	v%J-Q>��0 i7Z�j�R����\҇ќՒ�hO�>|���<��M��c�4B��Xj��	Yu��6���%��J��?���08_`QD���9j+�a��d���
ȀN[.d��OTvљ-`��o��p2X�u8	�^N�ve@�q�i�ri�%�1�H} �hցb/�6u���Rse��p��ć��v�I�E�@1�!G:	(�7zt?�i ��c�=�+/j$	�]����ʖ��gϑ)��n�796v��$b->I4����nGi�il�4N���WU�P�)]H)GW�;���'=K�HӤ9Dc˟յ��C��>����Q뙄IK��)pꑊ3m�����U#ʑ��!҆�(=V<���W,{���1u�#�+W��#ԭ#��T���@�S�s�*`���V�5�keB��{Zԕ�rK�kH�[�*��y{e{e],���p�v�)��v�ϑz�p�����a�a�Ȧ�-�T��RL�~�����C�0��P��`���<�9nd_����-��i|	@��	������{��04��~%(���W�@�m�^5���cq�� α��HF��9�sdtN��^2]q��gN �)_K����.RX�D�%C{����S��4�h+	o`���D �c.X�>lVFM����2�N+~���ч��|J�@���fE�������+����_���Q������s���^��p�������~���{%#���^篒�/u�����OL�T�9�{a��׾}XHs�L�j<[� ��-�"Ɂ$�%�GM�Ź�mp�l%�k\�г+$�.=���sF�o�q�i�����Y��[��
�����TM�����I���6�3m"���"�c&$'	�^d��D��W�R�^R�Q��$�
$�����|>k<����9��T��4Y�E�%����֠�4���.�l�Q چ�	P-���#�����\Zq��ow`8�l� X�$���|�ب@ι��^ތ�Y�\I^=� /)��C���c� �|~����p���+�dԺ��7w�<��x����8��k�␍/�Q9��i�zf�h�U��/�N��� �Ow�o�S�-����?V���:6��S���s9�`"�
��Ȧ�?��V@�\q������rG���l ��b��u�����b����!S{V��X(ן�ѾL����b!j�9�A������0��8r�{�j�Ѥ�NB�N:�$�u�%syv��
>��� �)����JF�ϖ)�!.�:>�8�f���� �}��TwA$(���?����~�]��q�h}�$���q~�T�>A�~ڐV��L����p�UR~�����w�c9�ȭ�'T �cH<t��2����q�d�@Y��2�b�n�ÆV�ъ9d�n���gCOha�AԾ~���t��2{�n¶�F��_%�*�J�o�O��.�I�gOG�	��i!lOc����x#b��A��_TF��E3�-kz�/��}���?�yTä�~_��72F5L�����z�=�J��XD���2�N�<ړ�;�F�0@ˤ��� �&g���!X�n��OT��W�6da��η�ߑ�h��a���ŭ��q�\�ӫy�U	bw�k�Nu�a�75��ٔ�DZ��x�D -}��ҭ�d,����d�Pa���?]]� ����[C>r1��1�
����~0sh�v_������BTۑ��$��|"İ�I�N<�Y�/�o�7���l_���!�#���E\��)��������f
�D��j���!����>�<q�A���uSX�ݦ��#��c��}�xCx)C��6����ዉ�����Ą��Ro� I��t�1w���[F*����������I�`T�
�G�E�t2QXr��,�(���^�L��*��,�z��N�B���k�˒���=����a�R�7u���+���H�N]�oI��Q.��N��
��Qs|��ۛ���J��l�s��g���\�@�'Mu3�h�Ê#�77IYx��&��
�0E
���ZT;��w��?�wS���XXz�:�H�UYNkm(Y+�
��.�3"a�TOd���'�~�۝�������J�u[�1����%/��1n,�v�V�;"n�z��}B��E,)-���u��rҎK2Kd7��R��A���=�x�N��T��8�Z���Ͷ��u[L���-N-*�J�XS0�Mo�C�*�$�+|櫖Y�g�S����]���Ni�r��n������%Z��wӒ��W�/�����#pWb��|�\��������w��Я������B��f'(|u�"S DN�3tz�X�`�����w��y{�o౦�N���Pw��Q�.���*��b��u��Ch}B��$��Bx����l��0c��@9��y;n.%	�OE�>��\���ˑ��S8�AZ:Tuv��p����5��1w�
�����Ƌl�(H�b_7Ҕn������&�;�u�H�V$�E���3�ڇge�rҁ.X��b�֢`k�]u*�@��N8WZ<��Җ�͔�Þ���C�1�I�I�u�OC'���ڼ;}�&�O����ԧ6����W2���/Ɲ�KMW6՚����NCv��@�I���ox:J0�|�`ȹ,fP �E��!a~_W_z���s��,r���w!�A{0�?��G�Г�o��g��Ͽn{���Ճ.LYG㸮�/��ˀ4��rř��-)�F���_�(z-��Z,8�uƮ|�eE5�XG�ɏ�M�K��-��|N�������Ssn��Λ�����e<��0@]����{��A	|�D�J�(�R��$Y���A�Q�N[�"m���󦁓�n� �l5O��VƯ仚��C�:ּ�oM�z�d���͵�Vr���jb�輩�Ob��F��&���%��,���Zi�yC&=b-
��NҝD#f��u���ڇ���k�t�c��N�}��8�Z"��ƚ�5�y�l�C�N���E��|����ޗ����T�����?s^�=;b-����0&�b���l��W�qP���q�&fuL���0egA�)�q�;���Z?���%s]A+/������rq���-U�C�4��&��#9��8����e�(��ۚ�=9n��$q.\�$�����Y�蔃O0��z�u��ތ�:/G��A�t:��������@;��I	�a������ed��YIۥ��{z�ss���ihİ�4E@O�w�AO�\U$"����K��I��M��T������[pF�g%<��>AX'��߉��X��fQ�s�}_MFґt�/-���
��\�e�~^9�����D��Q�����^Av���c�x�g�ΛU�-g?�s�4�3i��p{��r9�cg3ҧ�%�!e� ��Ibs���@�t�����#yL�İ46WR`f����Q~!�>U�@'����J��֒�[��M_��K�����5	��ᤛI�)�Ck�p�B��Q.$����ߚ�fe�&(U�o�������S�4��k���d��;�W���^~�7wt��6�l�K��qYWWX��u���Q�y���;S7x�{��������Y���<�w%熪f��&ߘ��P"���� RL���Q_U�T{F�Q��	�IE��շ'�n�#R�Q��{B4q;x��
��N���Ţ�]�Zh1y40"ֿ6&�]�D�U%.�X{��=m��*�k���Xp�#%f"��d۾�܆d}D Q�;kCGN��H',1������S|�ъb���A�A��*�C��o��\+�d���b�7)O�qJ�Y�|$���O�c�6��T��1C�{����1@x�������M��⋘�!��{5ڣ@��{_m[m��UK�bOTX9D^�@L9�ae9
��K?�O�ʟ�2$���D��	P��ORi+u��m2o�Y4�3��ߌ��ܯ��Q�̼˩m�t�;\脐����w�q��D�����?��8F�WX��{9ac�5[�	%"X#��^Z��BQ�
�7��{������4�]s���7<��+߾%	h�O�ZS[�ݠ�{�c�y�7��ew%6?�3�#�!RR��!�A�ӆ�J�&�>E1�iy~�����g������������5	�z�Z�#��n�`��������UW���Ӧ�|Of;A����{�`��4h87� ����4��"�k�k~���f�� �_���/Ә�E�y��ws��t\�O�Df�W�pmYJ*���T�ާ���83".l��<��v1*co9w��b���^{�9z��[�-��GQr�]��!�bWo��Tɽ�3S��EjhfM�2^$k�Ҽy��|Ж���\�.�ϊ�nN^����o��Κ��a���a"�C�����Ԩ�UΆ�4�5Hl�Z�O�$�-�٧�90�Ȁ*���WXU�E��&�~������_�+d�_i����~�>�toA��Va��#���h�!��{W+Tv`A�q��ih�V��M�A4�PH���O��fb�!Ϟ��).�Po�`����'����QL�"��w��Dc��ֆ�[&�:���V��ڹ�<�/J<ٿ'7�c�'��¾&����=)���`^p4s���<�JF�#l�IY���ÒY��0�N��ݵ*k�(��f&�m��"�m&>TM��\�v`�X�U�������aE�Mȧ��K4f���=Mp�C��.�1�C�����@V����V��_b��g�P> q\Х��`W����a�]��iC1A�wp>�^g�bo�A���"�gV4'TY��7�j;a�ȑ���#�9}��Tm���=A�ϼ,F86ٚ1Ȍ�,��C��=K�2C>�c��b�0Fi����j�3_�!�4C�=U\�Ch{���'{�+E^�e�MO���hh8�^ؤ��X�<r���∅&2b�R��:/C�4����<���c���B9OZ}OI	�)�����4ϋҭ��~�L֮�s?������%�	;6��sg�?X!���s(Z�f���ܢC^�������$ZE0z��3/lF͂�'ē�-�>w)��إ�����`�?���>e6*J��|~j<�9�(�`��3�y�Tż�5	���+�
�Ӝ_˜&�O���<�
<	@�p�����i\������������i���Bb�l�[�渭xk�E?ִX�=Y���ώr��������Z�Hɷ��s���>��?\}u@U�����Cꒂ���E:%�K��A@BJ�J#���tJ#)ҩt���>���?{fwg>S{f��"�]U�d���{J��ّ��ٵ���ϕ���^�a�{č(�H��u,��c�O>�i�Y�����;g���|���5��8y�@�.^r��.���5�y�9���冟Yi*c'֤���b��^,�C
D�J����k���\���:���ƭ:]μ�73oYeR8CkN��s6d�1Wfy��_�y�:d��Sq�}>;(O��eӶ���FQ6+�z�C��Do���r�l�\�~[EJШ��#]�P���<v��-���},QԒ�������?*�W}}N�7� �L��/�k���Ifa���r=�ߐ74]�+��%'���O:SF�v���"��� kƩ!
�<�����.�S�Y��z��&�'+s���/�~b�����W&�N�y���"��&1�t[\� ��{��g	'٦��Û5��ד-�@*�1��px�h5�Yޤ�ў���z+���$s*baR��|�B��<�Y&7.��E��y��WK��_�_��	+��������*���̹"U��m��)%�.y�7�.T��� [��|��@������J��+0�c�>�t�J2&rȳ�K���`mN�O��ҋ�<w��v��\_���J�
Pv����N�t8CZU��J�a����-�L������r:��#�, �˖ok��d t�����VdfSғ�*<f>���?c�"�rC��������{�[�%6��Zh��X��°�2��:�!�喯Z�(��+I�}> S�)k�.2s��L�c�1��ę	R�7���__J&o`&���o��+k�K��r��t&<|Z�����$v��GD���k��qf
:����^8}�U��m��jS���^�f�[@�� , zϙ6��Y�h������ֵ� ��H˖{������-ky)��,|���e^�|�Z_�%��ن}��o�	�XT����{�¨i�b�m�����q���\s?�ٱ�~K��*��1����q��x�Gd"FY�`����	�`��BT�]=F��7�'3����b�p!��b}G��];��m�B޻|/_�˰g�uq�!&%��wC�H���4�oVx�8���tnؐ�yx��y�5,���Y��M�z��Y���0S��T�b�������F?>A�u%���h^���nm~�v����R3���d���{�jp������� �,cQĪ��n��O1�.�E�#����~�6�}wfF����.1�;g&���y<���?����fSج����/V1�U:���.��G:X>������>�^oI���Mx{"�˾���Љ���=u�a�n}�(tALI��!|�w�s��<h�t|�;l]x���ru��<�f$�����ކ넋ll���z�J\�=�T�.����*�J��K�%U���fz��d��~�X�y��u-��g˅�kz�d}�ϭ6���w�s��T>]Rݬ�Ni_yH{������ɿOp=��G�Q�t��ryG[d\�n��>Kyu��,��)r��wl�n\p���J�fi�ތ��XՖ�-r�Đ��`L ���! AeߤБP��l��7��Lfi|�)AX��-Ҷ�g�L�8�ӣ|,�?/C3����Fp�O#P��H�ʢ��}eB���^ � L�L�� ��l��N	��5Nr���=��m"��s�Y7 >�\d�?ʶl�<ߩ�f��֩W3�	���]7�N֦u��&��@�(�Q���;�.�vV3~+���Z�i+� ��5��O��ܘf��bKXr:HI��BY��t����4z���T����˦'i�8�|�
�37aX����羬�R�7�a�}/H'��s�����О�J*�|����該��=�*��/l���I|O��ZQ|�L�ʅ�+��-�~Sv�Q�&g��H��)�}�sr?k�A<"�[��RBZk���>�N[�/	6">�X��Y�+$Z*�WJ*�T(��C�Ƽ���I������՞VgVm�/_��;����7��լ��g�����}�	���:�V��p�%䢟��K���_��'ۛn�bMJ���e]^b*��6�!��'	5\p��3|,-��dZA�S�GWp}�~���U�G�O%�2�����dd�bS�s\!bqqKq�:���m|��T����������-�,�_!�8v�\d��w�d�p��ҀO���D>w��5��
*6�c��օ7�>b#�����.����]n��[�V�m���!u_�`�.�%��#v�u����{��%�����54D!��DF�ؼ������ٝ��Q[�g���RRZs1���f�"��?=�F��VOP~�K8B�\�򎂪FR�ng�^!hSt.^&�p���~�����������Z�t��U7�*v���̾�f#�-����y�u6 �0]�n���K1q�����S���*����N��@>����HK~�������3��mpK���җa?K7��8��_����=�m�k_�A�2������X8��.�)|Wh��*r[�s@N.��V������.�hx��7=��k��G�1�D<V�y,?�f�b7���e���΄1�kv��ջ~�$�興:�P���R!��<�&��A�9Ӻ{�uZ�Vo}�"�;G	�NE��d�Xpy�5��o:�R�	x�wib*�Vp�d���na�V�(�.��j�O�L=d�qpR{��_�E�����*��˨< \��
Eq� �RBW�6��v�2r49E'n��}^/3(��CW���N8���T���#��l�0捍��	�ʬU�6�6��T���zE��fI��kA�sB06�rcB<��I��[���1�;�E���ḍcX�¶	4�8�~��RWy�4�}fJ�ź9��ơ��ݨZC>�h6�Yޟ��Z\?V�}��SǞ����\��~��" ������|��k�:���Ͼ�����w�=k�J�}^�4�NΕ��ϵ��g4�rwRJ�k݈[F۷:�<�WLR!-+X���Ǽzb��	�R}�u�/�9v�{�M	!J��ɦ�{�M�Y&Ɣ�b;A.a2�f�YTe�3сP�_Q�����h�����������=��e�ğp�B���6����L������Ul�3(fB �r�����I�jB�`i��f��C_k�d�^6��ui�=�h�ρ��Ѐ^�-�=��D0wNC!8�`R�bC�I*��� F�Iit�W0O��T���sW��+��'���m"h2ڼ�^o��l����D]�ÈMMpc�1�WDLe��7잌�8�tmF4xZ޴x��i��'��� ��Y-�!�\�^��!��D}�㙹����t�ݧ,e�5��A�=���xl� �R�{�$o��{V�q�,zt*o���7���ڔ�����ªz=�'6E>pDQ�1dS�����s�]N�׺��z!����L`��
�f����4-�)��sO��X5���X�t�VppЈ��7>��U���V��9I������sz�B���B�DS�r`+vm��"OmE����D�2#{hZ���k����TK�	������+Q����H�����x��􏮺/��j;�?�ʘ�b����U7�0W����&J������ZP'����=(������4>>-ٲ..�̘�0�M�&�%�c5F	K������c�̟�tӘ�E{Q³��	_�BS�y<锦��#��5���GgZ�|\��:��Ѻ9%� ���B���h�1���v���*�I��?�i��7y�N.�A����/؞zv<�)�<3a�f!n��syM6�͞�FK	�I�_rS�'N&�1�a0��OI�9��Ӆ����ヺjĿP��� �G�����|��]�)"�)Ȍ�E[���]�	_J�&H�\��D[?D��TA~�[F96���}��"M$��(n�dNqx�Q�i����+qK��W��h�܃��c�Vԍ[$�A��0�z3?p�\?�Zk�v5(�0%��6���U:i����&e�#� y�Ρ��D'WF��fI�!eb�����(����++�W+�ѼQ�������D���֓���p�cx�y65l w��Rk��f�L����]���?�M��K�E `5s%Ϗ��x+���E�&���~7�}Z�E���A���Fl_^�.V��8�)�^��Gɧ����W��&J�-YcL)A��=>�=b�������λ�K���oR�c�M46c�8�+!'�N���N��r����0Q�BS&���v_kF�E�;HBIFS�a�^���n���/��4���H��	qs]h�h���o�]����d@t������_�6N���C�G\���#i��H�Ӆ��,o����ʠ�E�t���G��Ե���� Q��Ս���� �N�ۍ�˦��qm���V$?��:�:gAE��6x�
?��}�7���ړHD�t��a��)�Ay�5�ݻPlp�����.�N�)0�|�2��y�%�i(��� 'ʕ��]y<F�2y:��j��Siʇkw�ǌ��a��Mw]Q>��$E-L�A�-CK��ZN&��$e��?G~~F!r�q�^�T�-~���̎�?07�`@�O,�L;H�6���:{�	�O�F�]Q2dV>��`�:����JWM�7S��*�U�N���`�{�?dG�ąl��b8t�ʭ`�)�tvZY��&�£]�S{/����U=�y�-�j}�׽���3A*�BN~9�)?w��ـ42���"9���.�8.n��ۖ^ XI3�\$���T��LΙ��*L��()v���r \�+�II��?��<�����;�-֠����pb֚��%6� ��CV#� �~�%f���X�b�{�����[������agp���D%�']�$x������K upϦ@Cv���u���h�:(���#�y�'7�|�XOZn�T����-��A�3�t��U�6۳��#Hp�o�&��(|�@��ӆ>sů��� �^�yZmJ�����k�$� Q�zt�g�:Q���=�_�pĦH��h^Bj�쪢J S�����{eb����S�i���*����i$x��Ł�Mz��k�cL����b���U���sj8����t*���%�`�>[�QOxĎohkK��3ڡ��yD���=bv1LF1���W�O9û�n"0.	�z)�c�U�u��v�-ı�����#~�BC�֛��7q�p�KRgt����-���G<-~WG��-:�oh��e�|��u�*{M"��qI��~V�3ad�iNDH�ɞd�Q�]}@�)a0��UI:q�;��9\�!5v��� �ֽ!ܕht`�388]�%�ʶ��@\|��e������(��!�����5H������X0�ڂ�%d�g��BvKt��|w���'�7YV7&Q���o�u{�I��Қ�@�!\;�B�Wkn54���ar���L^5=�t������C�l�9_CE�O��-1�ѪK��K�ڱ�T��n�]�z3�����*�~����v���PrE��e#�2�5.}R�Mm-���}_AaZ���.Y��������Y�Ve��SD��X�qQ�#���P�ј"~�?>F���^ #r�z��9�e��I0kYb'�:�7�)�dsE�w7&Į�,kp���s2��T��ŗ��'6ş��cU~.�"��I�S�b�**SB��G�Lt$H�;]���B�
Bˉ��v�>�r������R�iMB����۷ 	ׯ�2��t�F *"�I�!ܺ<�K� �"V� |
2�$��� �w�p��%�R���CMv�����J"jE�b�ď�?G1'�B�G{�0�G��#���*K��"�?���?T��6�?�M8�UH/~��59���57��Or?k��3>O6L���D���M�D�(u�(��:��fr�K:�!��V��8��R�G�]+,��i��5�3&�0Pp���<:u�1���+ }��|~y�� �j>kx�ӛ������U0���ЊɄ��&���al\�4ݰ��CƁlY�0K�����췳U��~��
���X�s�*0K�?��0�v��/M�d8��p�9�l��cjj��;��'H��ɾR#�Bh<,n�ҙ91y���s�U"���Z����GD��r��2��c�vSW���)�ΊD��:{�}c�R��F�����?�K�+�(rb�N!��a������3:[�LӾ^Ub���2訖=Qq�s�_���ya�k�N�i�/�<�?FQ�џX�N���
i�^�co����nyGA\�+#�C��K�F�7���gl�dA���cTAl�n��~5�BzB��6�"����1���ZJ�Q�V����L/�,T��ߤ_?�-�O�
�{��c�i*�\��Prv[EB�a{�ߚ!Pۭbq~�\q���w�B%�����8�A���fh��Vט��RF��Y��H��f�;�)"0f���栢������p��2�P�$�?7���C�o`@���&�B6]�<@Kc�xfI�x?�ц}}1�9U,	�$�<�u���u:>-.�L��ᣞ��|M:��1n8ls�b�<��-��R|����x����%�Jan��
�%Ww6��}�ѕ'��9���+Y�q~�:1'7���y�CH�.�`"�\�1��&`Ȩǣ*Ӻ����9���ݨ9Z�z�Q7@$�F�x����w҃��y��#��Q-�m�u~{��A�r�P�����%R��O@uafU{x|�q�5,�wqG��2l(����{/�	W^p����0l���}�Ml���e���9�5�0���X����t��]-�#z�4z�mw�L`;"w�לY[��Y� �;ZZ:%��J3[%	�����6ƕȊs�g.ފ��R;9/]t'���6�b����k�W�)�%A�}9n̃o�?P|Bi�Ơ������V�bT�-�c��WW��*����6t��3�o��IԨ��,3	嵝v�9�Y�^�^T�5�%;��Z��:��cR+p��YC2��)"R�%0�+>d�Lڥ*N&�H���
�؋�F�o��H�j+��<��7�i�͇�Ryq��,�T5������P��nIF	�_�!T�*�(U��n_,�ۥ�F�Pn(mC� �v���w�f�m�U�1��柋a�֩`�i7Ó�w^�}��=�a�i4��N/����k����!.=O`:HS����dE���m���F�0�&�Z=^w��y�����/rZ��(�7Z�M��=��Q�!ܟ��F�#�;<����gL���d�*�"�z#�g���)��E�^��|z��^�^�b��Q^̱P.�����J�ʋ���}ܻ�8��}�8��Ti�iG.����9<���Fpli����3X?���FY�aB:�����rz���!��lq��C�*e�f����e��Z�^�Xϴx11:�"$Sz�'� n��>O�*Hd��2l���<�q�<Ú+0G1RT{�-㋶z��EW-{������/Ԯ��.���blA�q{�K���S�$Ƀ�ϫu�  و�[m�io��\���Ĵ$��9��Mւ�`�$��XzM�mu���*����P�j�Y�aeBXX��b���yx�z�%%jY.���r��c�?�#�]�����-B �%�E�՗�T�<��Jxgk�
�M�L����SU�jܾ�Z� �������"�������9��4GSB7ߜA;��9�eͨ�BW˛��W92K��O��F�<���Y���cz|��?�$���Î�ý���c�]�(��i�A���}¢/a;9?藨հK��f.׸%j���3�}�F��~�� �<K�8%�B��'�7A�>��Ԥ��;��St\0wC.W��#��K�W�E��zއ�8��REq.��A�c�	���-��L<��xJ6H��]ۮU3TML�V{ź����3��f��K�0�ĔG���'���[.lR _L `���9��\�j�I��(����ӭ4)t���$q�@�a�	� ���n&��Њ~D�V��ݼ�v��e���^�e5~ݳ�~=�#t�	A�]�=	3���Cq�ى�w��7�ʻz�xD{�	��WG���nF�)F���G�L�7��\E]�p�,wG~����WL�g���ೋh"tI���N|��k���Cn��a15�P�2߰ Lτ����)�s���¼vߤ	�f7�7��+��1Y�Z˾V��𲲔���_����E��gS��P�7�l$(�Qq�|�O����� �����j`cљ�'+LO
�0�����i�8�h�sٽZ���S������|�:˧�A	��Db��hy㮅��rݗ��aj=�?�ԙ/��+IA����'6T7 i��qO�6{-�>�R�~7)�0���0��o,1��B�������\�!���#Xb��P���?Z�m���>�r��a�D?�B��x���I[1���3V�I̱�����L�&CW����8&B pW$P�r����&l�����1�)\����ѽ#!r��)�A�i�L4f���S<�MV��>ۆ}ht�V��U��	��!��zy���kS�nt�j{廰����i��a�RD[4� �'�kh�	{��Ź�/�!ʢ�<�5^��D.���@�Q��o�r��w9,�k2�\<�=�/�vIΡ�8��9��%*�������v�o�[���w�]��s��=�a_�N�G��2 ������9��.��f��S��紦��os*�>[L/�߸#��.���� ɠwݪ�A�h�g4�( ��G��
�9���I�A=�� ���\,��޲ �PV�|��D��d�_����|B�{]ks�ԟ�݄�L'�O��4�8���G�0F��zs�1��J�5"�!����҂<�_�>O+5[ǘ���{;��-�0��-"t��VDƈ��V�8,�vT��y�Df���-��z�M���K�/��k�@_����+~�|� ��[\�M��K��#F���c����j͹��1X�q_�k<�<R���%��(�&�����6�]��<+�*e�<eok�w�;��߼�Z&�H�ؤ������nW�o��KW��ܿ�j��Ĩ���@�J�i7��	簃+J�eל+�4��2��<�,�6�PYqb�1��P���	�pkB��ư��Ⱥ	k
v![���������	��NB�ѐ�ׂ�Qx�_ y�e�?H,��[s- �+l]Fc�q���/��s��(q����"��3��Q�/[t��Js��O��o~�>;�*�#}��pn�s������`�r�1܍��~	�S�������V���dO~Ò� )g�v�<��wm�[}Qv����=�E���-(��?�Ru�Xˋs~[:)u4��K"���2C�F��\��s�~��/�����	���A4��3?����8�Kwx���YN/�kl�i4Y��^p��;ia�ϥ_ �	�jҠ�G9�S�+��$e��!��۵1�h����W�C�/�&/L�͖�ʉf���q��{J0>DO�\�!+�% M����jZe���0g�`O�41��ym�T*x�kL��^��GL�s_Ȟ�������0D���^x��xk��g��#�Ñ���}cI��YN^�o2yn�E@�"K���������MM��-Od�C�A� "d�|W}�����-�W*�Q�r�� �<��.��]���Q�3�T�]au�zu��1�?s�x��0Ϳ��Lcb2X��)�gX�U�0s ~13R4�1�s��+ZĦm�e9���,�/�}��=mN<���#l*ڼI�,+�M�ٔ�h�4��g,Ѥ�5��}�y�G�i�qO���b�,���h���]r��. Sj�s3p�p/�Н�-۾{����m��7�8^������t,�oZ�e��kYP���R&6���n��9S�"��02
L�N�����kOi�e��J�U?Ȧ)��<��(
$)]�`��1D{Y,���pN�r�&lO��� �@(Ya�S'�*��1-�����|]@����=n6�riK�Ș�ڬvi+�D�m�҇�q)��&#�jvq�M�!�CN+�)bP+eN��fR���=��c�
<Ǚ����*���Grw��7��D�ќ�ww�z�P�пy!�{ӸM����*5TwH�*��iZ�#w;k�6}~'Ih�쏀�<r@NRfD�<;;!�_����?7�j�c�7����F��yۓ��/+xT�c�o�j����kZֆ�J
�k�_q��l�v=��G��͘m8`��������c�+��f7f��V=�˭E��FT�.��k��څ0�w��,����ߦ)������['�?�RV$��C��y�E�hR��h�8�$�m$�޳��a��1d�z�E�;�9j����D��H \U��m�{���v�G�����I��H";� �H�u&#7�v;�`g�ny�?��$��}��2:M�!������-�x0��HD��*/k�2�2������߻���F�h���M��
tJ0n$�W���B��w���D2�o��ҮF��?����Գ}\�\��^�8����QQ��;!��es��;��24b��XY��9�ϟ�9U';��� 8(�O���>���!��-�+:�m;a�W���\�$������oDRRgm=7:�]� ��*+a^5�Ad���IV�	�D�Jpt,��K(mԞM�^�ɂ�����}�(g��bnL3��g.��7�
������t�y�����CaV.T A�o䒼��T�a�~��:�Dl��%�Ǵ~�w�éc����C���x'�"�]�{m��f""O�
d]#�5\
�8��5�\\�+%=�y�m�fՇ[�[d����^2�X�tzr��S�w^�c�	����d,Ee>�lb���@?�|iD���>������W�O�E�b��-�yVA����}IJ��[��mz�����u=�WWNc���󵑔<�ئ�왧�Cz�A������zgU.,v�V�D���'�#�f��	E��h!5	ހ丩���C��XB����hd4�J?�����a�;'R�%iφJ���zB��-C3�M�p�����1X�9�e!H��v1���8��q����|Ko,�4����6ػ�����e�H��m �'��17�nCA\<�ҧ�����5~^3O��s]t�].��
nn�n��}U`IL�6=C?a�ᅘNLG�E��d0d`kDl�WE?��@�@�JO#꽵�ϱb`�~�M	�Pχ&�{�x��I��V
>�;GVn/�FD	LˠV^�v�q*"�߬P��R_8#٥\wiX�:;K�9=)����z���B�C��c�C���D�P~maΧ�Uy�_� ��K��Q8�j�r�����wB�,������X>�N�]�MLZ}�< �<�P����
J�>I��B�t�&[��%3����V��Nqѽ/��y2[���K���%��H��w[�'ٮ�H'W�jh����ﾼ����SUCcP�����m�W��hׅj��_�� q/�l=\�^�[�O��9!�{V�<=}���x9�Y&���p�>ۣ[�/2Fk֢^E�Э����Ah��Y@�L�O�e�t=�;��*����~\�$��C�y����Vxfc=U 5�~�� ���E;K��^������~�|ǧB��V����&�|�N����qτ�<w�̻���oj ?[o��T��X�=�G�ظ�S4��}6t����yL*j��a�OHl��|#8}��J����a#���#�lW��TK@��	*�f_�y��`����!ˋ"�h���r��Y��-��;$L�|g�>�f�t��q��Y.��ќe��5}�%�N�� -_�h�u!^��ׂ)˭��I>Y�7<�c}��|b�$!�8�(�*U��y�d�U,t��(ܣy1�q��9`�G��r�;s�����6��f���^�,a֐��k>�s'5)�n����\�]Dޟ!!ҩ����$�|���O0=��)[2��H�g	�����<t���@�Q�"*΀S!Ԥ�3�o�.�;W�F��#T�ue>AZ3%lW}�,K��t藦=���_��881ҡ�G;~D5q� ���?�職���Dy���Sk����Ib-�K45�d՟��_31i�?�;O<"�m����6a�Ju��e ���3Q��@`ɾ�}��M^��f�/�iw/2~����%��͌3��z���>vj�H�ʜcVw�g�S	�vu���V�&*q�����?J�K��CVbS3�Z�D�a�,#N�tj� �n{m9��g��������*��E��dr��y^��L���kWt���A0�/�G������m2�~��U����6*	\���&�#�7F3PB���L7G��O���q�~z0���S��>0������.5� �<|ztA?�Y��o	Ջ.��ݯ�䟤�5�\/�����ݿ��o�!�����=��_:W���վ�*�'��躿BT��j�k�'v�����kɲH���wF��y�$b��	%��ӄϕ�m.��h�������X ��Ϣ�Urg�0��w���L�g����g�P1�ޭM))�����y���m#���)�8w��ݳ��'}#fx/Sz�{�jba�BP�a5`K�2� �ˉ�\]�oa�C?:4��dYp�{�F�A��z��� *�c��}R�3l��u����"����Og���޹�{�*-K��~��^��3T�A%����Q]�7��2#���|�1\ؑ���O�u���&MK��1C̥]/Gp��Vio����zy�6Ņ���b�!�ý=Z���Q������=��N��%��"&^��X��w,)9��uF�R�T��C>��,|ks|�$e��Fw�CC$!i����ы��1;���f�ŧ_�����^����`'�����X.;��mh���TU���f�S��)���+�ǚqٓI���6|�Mk�)tGбx^��CP�#�nTҽu���'��&��4v�v�N�v��Ad�!��ax�ad�ad������D�m���*�A�/�נz)J�'�'��sf"��$�m���a@@<Jd�I���݋���^�P�}�ܳ�?�����/:m�;w	�m	;?��!���=Z�2JT�k�L_��K��;j��St�Y������mtL�fz�h��8I��N����OM����2�M�)��"���'���vH9�d�y+�7	��c_�G6q���.���3���fa$�7�Q�M�-���SZ��Ew�����jO�x�$Nb=(���?��,����ZΩ�'˂O"<�Y5�*cC(��mf�:�f�z9�Eve��L�W%����_�M&�6�U�fX�E��ms���k�[^�z(���u3��.��~��.�ɨ�!��������r�M+,V��7����O�#���o�CQo�z&4D��?y�t���b7\	���c��;�ja]c�T% !9
�eG*���`#o���W�{/��f�4�lm�*��-��������2D���*��]��y �g�a��R�b��Oc�|�_&�^K������ �KF$�iF}�јA�����Un#��u�"�&��ήV��'�O#a��'I��k��
�ۼR�c(E}�9�[n�~��m��ӺL5�,��+� P,�M���`����H�R�07>�8��x��Ѹ�� ��,̗B��oo�M|���j eiK𡹃���	�_u���[�u�>م}���I�[6��n��|��A�R��*2~�����?l����s��O��!��>�o�+uh�"�(�@S�Q�ͅ��ᓺ�K�1�#���������QB�$�J�����W��o�7�����no6���{����}���{�5h����d��4k�x�u����Hh��Px�id,(�i��?�i;)��9��A\v)����,7\*���S���<����)�9�����zv����[�5¸�ƮgɕG1�([��)W�^�"D1�%<�&����_��|B�Tu-���zBx���������T,8���V���C���,�8|w�TdL�D�5"�$��Z�*�B�z�&���.�w�Y��9#O(Aq�'�qf�e]�;���W�]:�	��?��#��_b��1Sʨ�Js�"�N��b����
aW����t��tw���r�'2��3_���=�ye�M�&����Q,C
=kyR�]|�u���ݢ�j�����<B�ǡ����lVua������5Y;<�EPC��πn��A��?��.nk��P_�a*�!��R?����
���0\cŷ��Y�5/lj�j�;�P�@���/���Z��&d����pꮟ����?}~KT��C�_}�w��lƝ�gV�J�h�{��r��نP1��p�Gq���/�V#%`$�`��겔���ߴ��*�ɻF�d�󳍍���u�2082��?\�"-S/�j�չ�+�t�ޥo�4\������j�w���
O�������
d,"�D*���3�2Ǟh���P�c��H��hڦ�ӈ�����!���v/�v�B߳r�(_��!�'���N��!����҂����i]V���ݛ��؈��Ki��>!�� ����J`��F��n�7�@��R]N�6]��a`1���BV"�T���U7���(QϽ\�e+� ��ِ�ֲ#��~�C�?���?�[�=���a��%")��1(qz�.��x	1zny�?o��}V+��K\M>k�h+V�I����pwW御�4���Ӣ�;1�
R�F�.X�vj����8�Y����㓄�b����������F�0��<�'��_+�Nw��K�oh�i�]~���;;��P;Y�n(^�9V�h��(�g���n^��~\��T}����7��wд�k�m�(��E\g��y��ܴvU�WI����/�<�<W����/�	��ӣ�����T�Ry8g0�G�'4ӟ���PQ�"~�+�OUz��hsC��� AU�/u�ڸu����F�*��������gO���o��C֜8|�*���T#~,(*�2u麇���8I�	0ή�*܈~]���dxg�(�TV��Gl���� ���u��fJ����@h������M���*Ù\<��A'�T����$/]Y�`�]*4��['�j�2:�>�z��ujp_����tf�gJ�p�3�������o�$��r4�ɨ a)���R���k�U���4�wު>��"n��-�~	V��S�5�{9�m�S��~n�����(����ȠqaIl�i!x�A|��>��Rpk'�� ��b��y�KI�Ͱ;�^�ji�g�9��}C�1?�IS����+�60@�ʖ:�(����rx1zӾ!�^(�w��ΧԸ��b��S@�pr����)�t�� K������3�Ԭz;o�OI'�{�3���妍�
�ӓ8CK��3�u>cʔ�s7:W��.ۯ4g)���%b�N6k��K��{N�������d~E��{��Ln:=%d��8[1=
K�ME����;	�_�Ǹh�ե��OP���'��A���ꦲ���4И��ث�O�>�a��0y_�d���0�e��9���!��}!�ST�/f�RU ��X�'�ͧ{J��/AG*�~�ŕ��!̲ٴ�L��V.,�N����`���� ���P���X��x�N�A�M�J���'��i_��}%��C���D��{Q���d��K��/Z���%؟�M��yex��5���.a��߲�~��$��6
������.��KS�G^��W�?�K�>�~���=��ۑ��a,�r����~2{���	_X�0�P��NA����	�1��8�O�g�4�_p�zJ��Ǔ�������Ԭ\��i?�bZ��S���K\E��U�n�L�擈�����x��=�H�M��\m�~���@~`��Õ�g�i�_�"�V�L�����r��m�����=)v�����H�q;Ӭ	�~
>�=A��57Τ����:�'o�1HU�-< Z%��z���%۾�Й�- BX�QY�їP/�K%�gj���O �I�`���g9�` R�x��A��"�L��{�	M��0��Tx����s΄=.Q�T+�f��P������F��w��ĶRZ��n>
Ǜ�G$<%�
��U?J����bT����(�isM��o��~��}���*��4L&� ��)f��#$/�]�H�s�}1���ӓ��y�9�x��6y�_5{D��'c�!�;�mb����nɖ����`��M���rM�]L�����<(Ȁ��1���������~����K�b��M��V��)���L�ȔDI�xG,+��8��>�N��4:���^I�Zo�G���T�Q\[p�5Ӟ|��>�����<)H�1h�?��t�P���^�V�)>>38�/�<���WV�z��"�V���ͫ�E�*y�xʀ3`?\��r�	?�#���ؘ�|�&�ql�0_��ȳ�)�͐3�=��\=�����f������'�5r�8�p*e��&���WM&3���n4�ƥ��=��EU]���:���i�3�Iy� �Z��7F�gH�	؏+��2�̾cbl�e?�%�hu�6���rA���6�5��."ؠ�/n�\���ٳ����y���ޏ~�e��m�f8^�����%W�uTI�
�2��|��d�W�7���Q#�B����W�vӉ����9��--�)�։ w�٦ݥ|�����&��S��*
�<r��4���,ɣ�+`J�7�	L�"��>�^�����r>ǵ.[�X���Ѝ�D��XJ��k4�Mo���˓��C�G��� ���վs���>맜��Ǎ��x�ݞ�gyx�G�<�;�k�>$fؗ���-�	>��G�������c��Qн��x�hx�n���z�[���祵?}4st"Gi^ƿ����>�Ęn�!<*�i���ѱ4�D����G]�EIJ�7�-���k�`��^�U�K#�t�
J�4J� (�݈ HHI(")��]C�
�%�3�0���=#���_n}����ٱ�Z�X�\/lY(��7�O�|�FZA.;�w��$��e�QwV�"�� ڑ����F'hL��u�TWU�{�s�+��qG-����t�g/AަJ�	�T|O��g:���Ay�,)�(�����ܿ���
HF୽��_E��p���R�j���O_R�OT���g��>���1g���ݜ�9�\�I�� �e�������-P5�!����s���R1�c{&�r2:M*�������2��h�����C~�?��&Z7��E�m��)��>>	OoU7���Fg��*U�/|���yn?	r���G ���c���/�Xј��zU�Ϭ�2��a]Ef��F^@��W��is�W��Miz�s+��lB�.����cSF�z%=n���CR�An�����[��nug����]X��F��dy�F3|����1�.B���1j�������nW�%Ⱦ�iZ�9�y��>�^_A���[������דe��V]H��X�t|��ZE��Kq�dp������iⅦ�,�)�!S�U��@�5��8�F�CT�m�r��,���,��?�b�gb�ˎ�.)D݃�l�_O�Y	��%WO�1�\��BD������f֊�Ņ�/�e���Ҵf +��O�4����k~�:D����Cʫ����W)�\*EU��\��D�j�&|�]���KMy�͔��m�{�1*��˗�e$��;]�qmU�alg3Uݱ��,~A��5�vp�����Q�e+_#�pc,�/Z5������5J}[M�<��y��x�OF��\6U(�:����E.�')VV{�K������M�S ��iva���!�o"G��@��YF��O\o��������nq!���P̐ʕ.��\4+ox-��(B�~;��˄�}` \U[����k�TEI��y��ˀ|������77�#pdJ'�Dͤx���K��ROFCYdFy��!c�I����\�PI�:A,bqٌ�ht]eM�'ϭq]I��٩\�q�Gj;\�՞��Jѻ�=?�"��+�����v�"���~yC���U G��=dK��.2�����1B��~D��{�U���'����,#!3�Ճ*�����rt�\Ԇ`ݻ� Zm#�@R�
�0[�_�?��J�.��Qj��e����A�:9(��db��]�u�<�-}iyp����&6�?b��YM�: +��G���wD/b�r�Ju�s~sͷ
�'�2oq���L�5��e��L}��F���8d������q?����.�#�����6�������Mu۹���_�>�f;��h} '5�y�*��*����������H��_������n��
����lw�w��7��	3��6��i}��k�2O�3e�u���N�����:����"m�vI ��Nu�7����w�s�L���)��C�V�PB��[^yr)˗X��zO�&Ȍ,��U,����p�z=��չ��NÞp�rd�i`-S9����^Ď���r�aVS�!s5��4�����,~����i��wK�eR`� ]���\��ت�^y�L�E�õ������ �z=-�z\��aP��iH�� �\�U�1���ׂ������S��S&��531��ĕ9���ޟ������z"�2���Mv���U��G���Ow�~U�Bۑ���4K��D�/|�hj�]������g���a�����/���a�}{�O[OI��g-��s{T���g�nʴ�y�Z��^�&:��ͱ�Q���+c���[z=!mw�𛿱1�-����T���&+�,"F�t�3���Z2odo4�j��F��ӄ�XxD�����p��͂�i�Wp��W��� �F6^)����c��w���	��$@��}�1(3��7Yf@m��trr��ڲO�+�/��ZrOW��H�r��?][��j��+;�q�y����g�E/saG����/��_L}�Q�Cit��c���S��T�����`!�4ѽ��}�l-���u�Y�pB���]8=��>|��a��ͥ����}��gH��1A�W��A,vֆGG ��<˞��l��6���т.�+��yջ���w�[� h�/�U����⫧sn�N�M�ʛ6R�ͻ93���߮H��z��_̿�2Jس]��`��s<d�sW��3������9Y��ֹ�M9�����L�ҋ�x��� �C���γ��]�����I���9��R���j�@ʗ�Fgǃ�J
33}��s�z
�����k��8�z?g777L�455O�p�3���"��I��)E���k��F���F�L !�`��@/�L��WUUV8�z���8�C�����#� ������$�Ȅ�@Y8�7�k�$��dS��p��[ �}���L��:�U@���%�� \�OL���Y-E�����\�ę�,��:�� H����7jr}�@�]��ۇ��>��!���&��f?]3.@+m�n-3�,���-�4\�[���B���&U�Lc`��"A��h'��JS�SE=�y��'A�:�T�?������~������s�X���>����Ʈg[�E48�Z��`���ÍWq��H��W�����`���x��V˕J�}�N�9�Mo�	��%Gx��)�ռ��(��3+`O��Ҫ���]M�Ϣ~��Z}�y�<&p5������/fT�0��ߣ�|��99�z\N����X�X�u�I�gx��2���_����z���]��8��<<c�*_��5���թ�`,�� ��~B��Y i+��[�b����@������}!�S�0=��h��D�)�0���׎��A�3|��SԵE~�<��_K<^�D^��`�����C��
���$;�fϚµ����}ĽN���K�.��g�$���6��V���q���s���t0�W��Q��g^�4�&��a���r���3��i��ڴ|�1��x"�64^X���m��ϐ&>`�j�=��x����jLC�WCz��Q�D�v1�-���ũ�kG���wvvN�:� � CZ ���fE�X��|#�3��X<�k[=�����k�ͧ_�D\�����?O��x8/�JN��0�N~�;�ڝ��[��ɣ��Eq��)-������8f��<@p�| H\QQ�@J`����@�l@�>	-o�� 1�i�H{��4�X�;��UYt��x퇀Q�K�9(6��������q�����;H�L��*�Xz��LMna!WsK��yFX�<6?L���E�����2I��T�!�@�y`d
T��:ո��kl��p)dɥ��M{/��f��[Vѓ��Ǆ�����jhX틭��~���y�~�+�T_,5/>V
3p�Ó�����rw3�z���m~Y"k��֝gg?��{A�k���wW'QF��!���W�+ͻ��Nm���ߺ'Ҍ~��)#Ԅ�52��~0��R����Ih{��X������x:�ڲt媤$�:�����PB�x+��KN��
Rͫl�.V2�GL���|´�9w�YA�m��@ʭ�D�����a�?\�[�2���?o$�5��l�>�)0n3��h?���:��.��o�(m��hw�)��P�G	@��~��^f/K&��8oc�b��=��V6F^� A��^���1 
@�[�/�uD��|���G&���g��K==����� oaa`�oS���8�Rt��?HO����3s�Jmߤ�`a&`ΐ159���mx����lfB�fMol���f�L�3��:�����:##��j��L3�O�3��TJ��G q��1eg�6��(�����t�K)���{8&Wmm�_/@�;D
��J{9��dq���ބ�[������v����?a�8n�qo+u�M��T�Bn�y ��o������un.Մ�5..�S-�jF=$止[|ǔKݻ�7:�i�5�@����Mc������������7H�O+�*��Y��ζn��:;O4�&�$�P弘PŢ�H^e5y.��(����g��s�,O�&m�pn�5�,.���s�3n���J�%[��R�2���kz~�شl�8��Ē��h֦�v��Cֺ���~�Z���KRc���N��Q�0�u�������v�U��^H�e-n�	�oxJ���^sm��rrTd����M�g���6Y�W��!��5c�����H:
8�q�b̈�3�1�<i�_�mEf[�-n�O����ɹ��f��� غ���y�
�A�*�����Z���H8�R�҆4`�3�v+!�8�M�|9���,�"P�W�Ld�ᒕk�\�10hZ21�r�X�)��/rq
|����h˰ޯ�´B�m/�����"�)���.�KY�;���G,#�N��V}wd�
����~ʂȝW�_�FX��G9ۿ{�I�RGD�Q�A���X_�r�$�̥ԫlJY����|�r|p�Q?�hU��u��C�i\򳑫��*�L�!?h�U\�O���m,,sm��q���J��E����ҾK��Its�#����lW/��1�8�������?P�y���M�2]-��s�nӬ7���>�̽W�gNa�/O9���m]ʠ����������%ޤ��z�;� �ޅ��Y��v�+�G�I[
<�b19(ʴ�nwC�m�R�c�'C�;D#���3J��B�cY|��o�ʋS��f��ϛ������3y-�OieE>��L$�юz~�{aO�*h^���-�r8�+K��0g\g�|A ��/�� ��K7�� � �>���mh�b���� ����x.��E#�k�>CR��t0ا��Sʮ�`F'q�-��?El��R[�>��]�*��΍~�d�[�	C��x"B>���,�����6��H
GI�5���O��}*~���<�q���#�[�,9q�r�K�nd|������@�����K]?l%���R�Z�*'�*�^f=�����5���)Y^����?�\k��߷��T9��q���P�:O߂��d���"9s��?)Z�~B�Uvϟ�N�6��	�&��2�w���v�r�/��*�9�X#�&r=Th.l��8D�,]�d���y6X�֢�Gu��T�ȁ�H� ��ʯ�p�"���)�Y�^�j�^�.j���st��o�	De���S�������4�mVr�.�B4������N.�=�Uu�ߛ�����k�`�6��? ��uD�P�j���B�em��.�T�3b�ghIRjv��n00�
��wH#��i��s �Q�j?k��%�V�(�����#Qtm��ǝE�W-�4��JETĎ�ϼ���Vg�Y1ί_G@����Yml#^9e�3oT�c�
2�Ł,�����J;9�3�hE�] 9wO�~���f�*s�b������<�W�����ͦ���~��

�d5V�E�iv�hme%�	fP�"pe�|��gqŶu�E���>��Q]E�$����Gn��BaV��� ��R�6���ry"b�%�yl �P�t�-/sD�:;۽"7�ZX����Yj�k1�����4*�T"M��P�wZ� K�b�\�j]��!aΈ�ð�Ŕ�*��a?������~<<_rdPN���K+d��"X���Om��-��?9���ӹǛ%(We��9;Q/����DR^�Ŗo�*�i}5�U����|��H��o~�P>��5r��j���X�`�gzX�X����{?�����#���w�J���h������z�c��}�n�{\s�B�t&�Cs:����j�3�'i���)dA�o|�0����GDaM�'�>R���l�M��̉�[^�j��8#M:9�T�����P�Dٝ�>����#����{�!0?�bv:z���(��3p���X�kR��E��ww0w���G0ݠ���z?c�|냜q1�h 4�66T���#Ng�A��l	�u�ϒ���>��`䂆/'�%����t�k�����3�=�ޅd�=��4׸>���6kP��
��}�y�n�g�g���0w�0�{�}�I
�����XX[J��J|i�c�=�SI�O�ђD����^��k$`o%i���'�<�(*-_W��K��� y��aE�������9�?'[��NF�$�A�J��*eB� K��x%�>�y���msP|:yǁ��૥��f)1��>�~�c�i�^�ت&���	ϫg�Az)�v-�@��T�Ydz���<C� IFW�[��䠵R�%���\����i��߭I�/7a��PH|����]���g;J��T6�t�O�n'��"��/E����>�Xճ%'r�i|7�|��_Y4���PT�%nc��
���S>,�C챩bM�L������@Õ}�eM�/�i>��%�$ �3}�#��o�m$5�����<9��9ڱΞ���S��M��^��]����*,%i��vs ���~g,  9�����f�b�b	{�٫�"�E,b����[�R� :U�ٺ�疯o�9�H�����N�S!�T�w�����W���>&����w|��Sd��Ծ8��Mc��l-
��
� �%2�WY�ygb�T#*�0��l�{8�G`��H̑���3$����
`��2�<���z*�+� 䂓 P��ް/?��btJ2�	������.�"�ڀ�bҬ(��4�m��F��d3�Cy?�j�NF�f��O��Q-ЛZ�}B�#��L���޼
�5�i#n}�҆�:�CښPh���ȣ�L�|\��:��(�Jv�[Z���g��v��)c:xiy�,>��<6�W�P�$Gp�B�(Uu���/�ǧ�XOe׸�af�O��6������k.
��}
Ծa�\=�pL*�����=1W:������$D�ʣ/lxr��nk�����'�yhs/O
]�[��ޭȤ�E�Pw��i�}�/�1��_�0��0�U>{��@V�8�l:�s��M��?<���H��B'w��&3��HĢ�w:�m2�t��u����L�Ibn��3[�gKy�����:9H�%@� �Mo�/9�s�L-Q��ܙ�T�J�=J���8�}�}��T�����'_H�Iu�RB�����}>4� ���D+pG'�2�	��yR� hQ�������x�g�I��#؈j�` o�����y�4�,w��������Uin��� �1{����"��/��%�@f��|�_�N�҃�;��g��|�G>�8>���C,�����7����\�S�	��Qi^v�[�ۯ|��lu��,��n'N��T����f��f���_�SaIĢG��ʖܑ�I��#�������SG��^�]r?��|��}�{�
]�����s�z��%(��/Z�ο�mݴl�JӮ��y,BZM�|�����k�����O~Y�}�ĥ|���E���ј"->�Ҧ�m��)l���,���?7#b����]��'�h}�~���{AqmNB�x�_bҤ*O��?�Lp����NV�}_�{�(����r��dȜ��џU$�gvg�nڏq�Ѿ�퓲���xji��u���	qYA ��3���X�����;��^Q��>� 	:h��Y�Q���Q3��b���Ё��NI�rIx;�EX��g���+�0v��~���}���,�5CL�;���?[ �Ҧ�m9�>��8�A핞�7N�oR����z� FXK\f4[���l��u5��3�T2n�c1�!������įDwE��Y6�"!h��-<q����#9��{�j��Z���$t����!��օճv_*}Y����'M��X�L��WS�����
kB�A1�7H����9:6�bW�<�o"h��CN6_�y�=ZH�k"��vG��R��v8�]W\;z�Z�U��ǩ��7��&Χ�'J�$��\�\z2Z����6�+���L��G���6��f��C�DY��R�?{��,r
�`K��a,�V��b"�S	?��+�-�+k�� [3ȸ���������,[���u�7rЗ�8|V�����{���r�o����W��Y͜���X2�����%�uG&i)ԙ���B���R	>�|��4e�T]�B4w�q 9��lX
KL��G���
_���e�r�8'tU�Hye�o�ZDWz��h��v ֑x����	��>�i�X�@#��&�J�+K���r���a�<#����J Z��Z��JX�k�*�}�&������dnr`��;K�52���ƺ):���˛|��.LuJ��u�Uz#�M��=�cڹR���L�Tx-�O�~���|#; KA�"?��
��^L���3��L�f`�]dy�L{�M
6��v$��H`��BE�f������H.T��L��ݚ��c�奨Xp����.1ќ-�l#�	DX[�_�w%�K��"��|s20�~I�(m��v���������h�����^!#2�*Y�V� #�3���H������c<~���	��Ġep�)/DKRr����Y
k �=+J�J�t���[�h.wH{������	ͮ�e!����-�U�L��Ż�ݞ kP�eޚ��fYe��.�"���O��XFv�����L7�A�lC\����H�����-��O��+Me�� ����rN�g�¤��N�;��$o�˚`�R�Tʎ\��:�����iO�}�w��+Ow\�T^�D8r��֬�9�_�u��Ӵ��p� ����ך�]�Ybs�H��s��U����~���lg,q�ʣeZ�%}��W�1a[+Z�A���Z����)���f��iQ�R˻��v��'*���r,ؤo�5�Z������k;"M��X��e�U0K1�>��|HNĬ�3�^G�3��[�5��1��ŉOP��e�}���7��5~X�lI�3�Y����X��$ʡ��]s��la��`���W�d�0���&"w�Mv�wI��p;a��+��1�����97�s�iu'!�Y ����.ñS��������fQ��	+H(�O:�?�Ӱ���B{���]. 9?�y�!L�l��jK�pɗ%�P@���������6���KU6�s�?���,��9+]qi�]v7��Z6H�|��ǔZEz�S��jI������t�cRrԚ���|Ź�X��܀�h������*d+��Z��ʾ�(F`T���69�j��t\�A�!�E��T�[���'-T��\D�t���-/�&@9�̴`�^��V+���R�� �����Q���ƖP�?��b0��əb��;E����#
��Q9�G�e���O�K!-W�)�6L��%����������|+w�N����Jg�A�R	k}�}�hۃ!1
��b�,����O�sdE-O	Z9��h`�����Y��3b N:t�{����"&��j�78�[9~�_�o]� iG}��#�(�k�Y.^�%6��)��o�����fM��_����'����6����
�7�� ی)���"��K@�CSS3+�`ϕ;y�����k8��~կ�-��ꝊŅX��u&�˃�e�6�~�*`|�B�΋'���,�g���z"�v�X�$�O,�m���
s���pڏM�W7��ar�Aؠ������U�"����p5�bz�.�����"��r%XݮEK��-s��Ӯ�g���C?&�D��V�|!c����b�UP����I���f|h�孵1�����y񋸫�;��fM8��O�5�7Q&<�O��$%�;�z=Q�ez�p
���Q:.� ��:U;+	�Km=)D��9^�Q$����۹�Kr�8�	k�S��t��5�md�&�z��A��;�5�(TҳP$	�`#�6�J�n$�y�R�4|
�j���e$�8p����TQ�淌�?��D4��fw�޽TKV��|&�O�&9n߂eXO����$Uw��Pi_�T(�Ҿx�葖N8�[�}r�,����q����x�y��hA6���dЍ�_ћ�%WXe�'�����5��c��P��f�A�#RAR�L
�&
��#�(8x��Kم�J� 
��tk���(Op/W�11�j�g1���9�y�����Ac`�G���k8Z������ɂ�g
/��F�Y�������X0B6E�*ƣ��l�#�A��N�oY;W�cNn<Q��_m<%s�f7*z�T�3*��b8�SQ�o�A����.+SZJ���$�{�]i"�ͺ� �Xw�C�gF4Y��L�R�B�?��Pз��ի�Q�����"9x�.���;�����Eę�R�;���xM�v���@^�Z%Eg���\@"�scij����A�����]n�\�R˃�HE�,֙�;��Wޞ�sA�t�<�{��t�vh�[`]cu�����0$��w2p���_r"���~�3��@�A�8(��T N��-�7�v�>o��=�ZD�9@����H��?�r�J�p��c��b��Ə����������m�V�@�%:saz/�?��v��,�e����=O��ҾY�E�8�2������:��ވ�1����e;�<�&�]��k�g�j6k��o�Ȼ=Z��[�����ԫ(A1&�6Yv��_~���q��(q	����zl�/m�.b�'C��Ǯs�h��R���h.����+2��ߏ�<N�姈u6;����(Yc����)�dY������X�$��??��� �c%����Y$K�·Q�����0�y�}�y֞����l����+.8�G��حd3̎�aa{Xق�Qk����H��v���&��!�lK�h�7?ή������������ſC�G�܁�2I��H��h�pC 7��+��u�a�6xX��x2�m'Z���WC�O�H�V6�����z��@�)���������<�i ��9t�"c�zO|��-oVE΃v&^�|{�c������f7؜
����?8�տ|�o�
ؽ+c+61��l���{Q��$�l��Z�g�,B Y+=�X�N�a�>�x�TZ#w�2*�@����b�S�o'"V�{>S�������Q�ءZ!�9@w����x�*'�}�aMV}Y���8]6!���ŗ/��X����`�������]%��K�1�T�E 2r+���]Β�a�Є�x�]?�8*Dȥ�cw��
�J���X*�k�� �OE�wr`[�a���FE�Wx�g���5��FX(&Mw�r�&���t�
�?B�4��o8/���e�@�d�|��'���Rf� ����
JT��X�L.#6[���=���=�_�ìv�R���}IX�� 
)G`:0��/+a����\鷈�R���y��D�@Q�81�n�_N�cp�g{,d�Zᩐ�>Q�+	���C�;f��~�-#ώ?xN���} _�˱R�~`��:�7��bFg�v�B��
f��'Cᑦk1�k>�!�v|x�l(�T'���Q�L����N�����*��d�xq��ɿ+����U�1F�\��m~�P�=�ڗ�?��w+ "�ޓ�����R��"�j*K�[@���#�^afgXΛ�Lb��h^ܰf��� r����R�&"_��a����)��JGk�&��d��g��u�I����@�r|nRa�@e Wu",�k�������$O^�ڮ���Û�u�Y&&Y��I@���b;���c�R�h��y��>�~�P��2��v[�Td����ѷ2#�M�*
���P�����UϗY�kʛ�k��8��u�{m�~$g�r��T`g�ѭI.�@��_��'�Iz̼#$�@:�5J���/)i�Q�e�.�司{�s��<:��XN�� -�߬����$o���M����mN����~S���'�&H�{$����pG���x.a�DI�F SbN��{uy�C#�Ng��dJ����3ɂ^�.JݰEv,,�b�<}NTjֿ[a_`�%,���&�3�:�����*�Y���@�_�i�ݺ�&sN#�1"����kq����H�&�mA��Z;�vU?���}�>(K�ڻ,M6i�����iKߐw��e�,`��i�|���1�F051} 7�g z�?O{E�����M��]������r���͘ҹ�~�9�H(l��2q��8��|��������@�t�g"S�dm���Gз�r�w�z�X��*�q�v�/�#��%Ȼ���L�Q�v�>֧������ t��c,.�gA�}Ȏx�ލ�uJ�{�W��U��a��/��W���$td:?��#��:e��1f�r��ؑ#�u[�GK����v�*�d�Ĕ)I�B�>W|p�/2:.W�{�u��2��8�H���v���:��-H��B��������I����x�(!�
:LA��z�>��<�e���&�s��������� �l�a�'nM�ܬj�W�5�	�	@B�Bz~��;��C#�8�J��YD[�*�W$���������0\�ή�m�#
Qd'���P��t�[K��_)�N�%�1��O�PZ��� HsEQ�#��'|ҳ�t�����u�@����t�[[�F�M��;�(�:y����Ԃh�S��KS��������Lj��[s�+/ ��"����5"� �n��\4�?_���hԑ��2�+�WMW��wW��;�yk�aRz�y�%W�t}�F�n4?�PT'�a��k�*�E����j�'�O�I�!1��@�xeQ~�Y���&FR�P�ϓ�cC���]�')������������!�5���c�5\���y(�k{��;$�NCl��u����#�Жp��dA��0>m���#�ۿ�D(����R�	l�bIZ�Y�?��h��l�מ��N�F�S�w�!P��sgλ���I�������
z��P����������B���[��$�*��RfOo�$vO4s�d�{��[�L���}R>�X�����{!��k�{�#��4�Y���Y���/���eVs�"��⣧�P�u�bs[��͇��j��Gn���#��DC��y���!�y�aH����hJ�L�r�h�1u��,r8K�UD���!�)�w��X����l��B>��1�u+A��D����N�$���Φ�3���bSt�x�p)�z:G�;7_�䋫�i�}�J��=�WV��ڣa��5!�Q�7R�Y���JX���S���Vux��-B�n�L)�.?'lՐ����XQo��ЩRߙ��p�/`���3܂)lPp��	4����q�S��L�
�/�T���O�.��P��Gʂ���
(�]�ϹO_*f����F)���Johԯ����xb��n!w`A�N�R�XlX��F|��5u��:X@��E*���0E�U�$�T[��>o�ԝC�	���_�� fN��r:=�ƎrWГ�(*:�V�~�ϱ�Z�T5�T�
��~q&I���ؿ�a�M�ޚ	 �(�������?�+k�B��<���jG9z���]�'4�:�e�$�ⶱ+FwT������$�-d*#��D�X�R)!��C��rC��I/h ��;*�f�ۨἙ@��Zfr-˶zFH�H������S�P�4�}�xc��[@��:fg�zU�-�爏��P�&}崼3N]���y&ҭӷ�i�?F],_0��Q]�o�؍�/5x!b�u���S�ς���׎fOE$.�?��~�]�ӑ�߯[/�S>-I |l�����_j���pͲ� ��4���#�T��3.�9�9_��@�/�i��{x2:�5���p���c z���Ѕ�l{^7,4���z�v��J�in*y�A�ǈl��d����֕�}i���㍆ϐU�
*{��z��`iK9
�m�o�Z�ą�fs�W����E��������x����S
�yһSV[)S:�M� =$����<���L���Z�r���dg��b(�U����ڞ��٭ܝ_yo+��b|(�ܛ�QUfu�������JN�`�gqFm���Jzv�7��n}���K-4X�Z��6c>0+64���Ҍ~Y!��s�tb�	�L���#�y7�(wD�y�8���sYLy��+�J+r�.2io�
��-\n�h�i����T����M���*��+Q�Að�WP�V��&�si؋6�3�AbrTRbFlGE˫�-�s*<�z�)g;L��Mv\؛�ARP"�	�{�,?��v�>�ɶ
g����y�;$G9�r�����D�'\��ә�Uz��L!����r?Z��;,Cs�.�q�Q���ۊs���
?~���A�}]�F�y\)����L�٭�����B@?�^����w�t$L�Iu#�����������0�������
Je���8�8��$�N`���D��Ū�å��K.�w/�T{��K/�S��&^�\_��圿:M�8��ԩ
.�j5c<���7��,���ދs�ro��7��3<���]�' ������dCb�&}�R�۩`�?�HKP��x�A*"��HS��Ty_��o��8xw1/�p9��M&}\Lj����{
�m�Q�l��,��A�C�\��ᗈ/�Q��	��<������T���e�Y���6N�d`<��u˼�i�~�����b�l��2l8�����PTb���քxk0���LSsarS���Y|Bk�W�a>��F�|w��� 1���qS������߭ZG��G�F-U0�V��Ń�l���ùX��K�Ҵ��Eq%V:���jߧ����+>�@���{���IϤ;N�_��G?��x��ԟm�NJf��I<�� 5˯�e�~���������>�;�?��I�q�����H�"J_�Ł��vގ��ſ~�r���X"����w�0������ºe^�A9Uݲ�a�w9�Q�K�br~jD�~�Q����v\��d�˪���t�F}��+�c��\�|)�Ŷ���f����|�����Q8�TO"���I|�p�<��G����H�E
:&���&��?�^U8�O�z^�9>�>M��Nv�u�e�=K��(SH���5d�p:6_�v i�O^���X,A�baIj�b�g�?���ө�<'t��L�H/K��(��' :E����7v%�+��ܘunPYr�~6kq�ᢿIݷb��{vj�>�6���Xllw�A��� �m쎠��GM_'��?�_?���{]g_������+	�u���0����	$�zSiA�	��X�`�sYX+�ǯs�Ϥ~ w��a^��<�I�%�p��7��Yi#MS��$k��ޗ��5���?�����n;a2�111qc���#9s(���;;��%f]jW ���ܥ����e�|����>�f��]�S�Į���N8>*�����y��4��>2�I3�Q~O)P+.�P����%
�E?����ӵ�"� ߗ�,��g~N�uq,D�?'�m�Tnl3Y5G'��o].�j����w�b.G�fҖ�����çm@���P������ӡ��{N@��[eMM�Bڎ^�,��3����]���·e*|�s^#e^�m(e����"���"]T_wz�4[�L�܁���߈+D�<#���x�H9�4��:���$|����ݳ�Ҹ�<��o3O��K�E�ۍ1[f��g��Z�&oTnϸ<�T��cU���N�W�x���J���8V
'בQb<nV7c��lfKLm��{Ă��F��V���'�͞��W�O�oI�Rԓn�$��5���ӞFY�>��	��y2��d5c����b=��s�]E��e���������byY屮a�4���6P��%ft =�){b *�_��:{�⭣]����U�C^�͇��$=r�Ҋ�8ïKvCr���{�c�>oɔX���n�U]�ý;+�m@J�5k,D�N>uylJM�O�칹a��,omÑm�����Ny��J��K����y���`�`�.�埽\D�+t1��A�Et���rp%?��l��Eb��/�n���tT2�-���`5�^A��S)'��V�"�)�;�h,�İ/��6N �7.�,!��,n���GF�)�&��>��W��t����';�A~�}��o�Q�ƽ��3����D0�W.�ADBr� Q��r��aQßƳA�J_���`D�Bۙ��ჲ ?ηo��%�3'�?	%%G9��q���=�Hăf�#Tߺ068b�[I��n�#��	�\�D'.�9X$��cݸG�p�����(:vsʞ���y!�*m,:���z�=�A�V�f�FR(i�q��o�t�6������,����PU�֗�ϐ@A<~~�S=&`9?��_���^Qn"p���h-RD͑A�����Y��c�4�kק���oA��;��E��f|q�0�i�!���6����?�h�I�Kе����[���6��X�6���%g�r�Pv��j�^B���C����@�R��B[+N����3�n��J� �:�%��ӭ���oor������B�c�Rs���0N�V*� k��^�za��v����D�t�>��	�9N�,`���K� �&�$���5G��hH�#���'K��2�����@��3+P�p���y�e����(v,��o�_���¾���r+��/��X1W�#j��j�>��k�-Q��)��1�N�y�aA_���:�m�>���׭(b�B�E�ܰs�9����W���n�=���n�V�lg��!��yeq0�����hrZs���_b��ba-�guJ�wF�Pq��W�r`Ǫ�FB�(��������<��g���� ���dU$����c������u��;��u��JR��M�w�fCA�]�2�B:hӼ��V���g�N��2C!�S6��R��rz�݇�6/��L��s^�
T:�t��q�TC�/����4�8�ɷ�#	�{ycY�L�ܴʵ���B�o%=�x����y�a�_�gVz�	{��Jq�&��76%Au��Γe�f��*y��+J����ޛ�C�v��/�R��"k�v$!�v�J��mT��'�蝢��(E��}�d�:�Pc�f�f,�;�K����������������s�s��s�s��^���_���J�����I��ƴ�:z�U����7�����q���!m0D��ݮ�蒖��c�m+����-��7+��1�+u[/R"���7?J��9����������r�L7YU���iV3��(9
{���eK4	ӑ;�j[�@���gÖ��}����Ӛ�E�]j����Ұ���<�-<��w�p'�$���	���cac#c���x)ϣv5+�O]jf�X4N;0�8���29�۲���ڰᤥ�y�,%�S7<��M�xX6��s�1ګ|������I��שּ������W�����ː�&��r�]#^FIjGc���s
����uι��׿�Ե���Xf�����s�d4wE��g����U���1�����~�~�yc�9�W���skKNn���2c�pu%�c1�N�HA��s?o��c��3�*�m�z�ޕd�3�,��#�n���>��[��[��b8?z��3�ĉ\w������_l�.f<O�g���B�/|���M��۩���췍������ٺD�ܗ!	�{j� �ӫ6�Q�NML�9�_�Wr�*�f�is�I�����]��D�U[qf2h7��c�"���@��J:>yCx�`����9�/����.�w��pS`�>�G����`b�C'6�W���;�^�E�Z-VY̭�w��JF	=���9��\�`�]���'��5έZ�~A�����_�T�|��o���˿�[9��f��+�T.�M�y�^���%�mj:�����cOC=*�<4hǚ3���b�K������������ ��g�W?�ѬΝZZ��(�)����"�o�-K�W_G���b�鷞�O-�>%��n_O.��y��.�ѝ5}=+u�y^�/s;�d���˸ysv�Ȝ�7G�G�W���S/�d
b�����oR|��Zj�m��9���+��:|�Q:-7����_H�-lq��~]�ċ�W�_y$e�L�ڜ�Q\�Fx�=J}z�zۅ��� c��Su'
5����7_�q/������>/�� �
�L~�O��V|/��I�umEՎq�1Z���|;kM/Znuk_ؘ��R���Tt��|���<a/LF=g�����0ۻw^�1��>���mҾMR;�ʙ���q�C��Y�22�a�̤ꋓ2����Եl�]U�X���=Mʜ�EnSq-%�Ѷ���%�_�yP��~p�h-�zF���
�Lb��N��	|�n��^�l×xb_�I��;���خGR��_;��m�2կ�%,f�i���{����ޭ��n�������օ6��cY��2L&J��!�}���i<8T�M�΋<ZDiu�$�Jo�k�)`�._����ܥ;l�n�OK[��)�O7��X�g�����D�c%
��Ԕ�{
Wg���UZ�՞�zc���W#{�9�ch�������?��s��L�֙z����C�����<�ff��u~������|�$Ffc �hڴ/�u����P�z�&֟�m(���)��9ɛ�ǧ�Ǉ�J7*S�+ޅ݋�h�­��g���Ͻ�e{�BOY:^�%�D�4Pƽ��N��}�1_��r޴�X����E���*�u�D���&_,�w%s2F�G�:�:�ޏ�V�H�+髟�[5��>|e���dw�Aj��)�8�[�|�O����~�����,+~�7Q$���/0�
Ͷvb0Z�F��cV�ݯ������ӭ�~��Ԉ?�on��B}��i�d\�r�s�q�}�E%�i����4��Gj����W]���[Bw�����b����D8�a!��5�v��w�V�#��hˀ���}:.Ǘ���Ɔ^U���4�J�}˽�.��)�y\�@�\����p�(F�1ổό�ֿ�e>V>0����4��묤�y��d������O�υ�=
�>q���zR�5��nP��zV��۝h7���S	�}�KD�)�ǧN��#.\4DT������;�m���|[�@�O��f�ǋ
�{S������?�A��xr�u�I���~��Ĩ8�����p�۾�z��и�b�X��l-|�}T�Jyf�\�(��[�"v�R�vD>�~I�H���x�k�<�$�PT�kB{\M���B�]�N{�9]5oiRR���YY?�a>^#���QL^�N�'M[�E]���:�:�g�����6^oZ�r�y�'b��aY��s�.�X4�,}���ihbK��w��y+��n|�>ʵe#�ofO���&�a��ΰ{��>h �L�>�>	E�w���n�9���6{�
�o�3�x�L.��wv����7GDb�]�z�a��n�h��3-���΄x���.�/�ʳ��jVa[X�.�<�,&�q�	����M�s�{���s�aq��a���}Q�O*6	��n`���T�d��5 ���WeW�
�	�<��{�����ۻ���g��Q�y��p�������[��[��7�3�G�_��Q�*��;�P��_���z�s��g�C��E)Z�Q�o8�J��eS~�Z1��o�Ck��n�NML�ۅ��v��]�d�_y;��6�SnI�A��7J��K�Cj��1��sԖ�|.��Yb�y5�"߃��__�ל������O��Ӊ�R�#�E��Ϋ�ʧ�������i�ī��e܎7�b��Mc�h�����myg�6�7��hR�D�,l�^�����S�l"��j�_�ϳ+����&xwj�g�v����ô?am(�`��	�]�񦀐�}������ߺ݇
]�M�����ɠ�h���g��O�8��+�?s�z�ݪ��9�ߪE\��w)��9c�7�0��ϟP	�O_�i��ƣK$o'^xh�S���P�zN֮�|o��.̒ߥxw��y�\�%d�i�H��/و��G����g�6?6�b�.SYO'����wj����+r���=�<�홱�K�-�Q�O���s8Ɍ����Q�cKʳ`�Nx$�g����������U��#c6�������ʡ[����v�K{L��)��Mt=���܆����$���ك0Ҫ�����j�ɟ\�;+s�b�SG/
�,��mU���V`Wf�������>_�x���iv�.���_{�V��Hm�K>����j�qS�����+冋�4t��t+�Ժed:�w��hy!g�'l��JÎ��.v|���wb�/N��11�q֊����=�Q�6��o�vM������ҷ{������&q��^q�iDA�8a^��>�������և�*W���I�T��k袘��Ч�,l������Rڷ9����i�&����wO�ND}r�{>g�9z�i���b��D|Xe��J�7�=:��/jlx��!y�x���r���=�7�YR����/(�������������\��ϧ'�vPW�����=ee�t�x����i�~�-&��&��(��/�p������ZZ���9���a؋�k�Ԣ��͙뿽��4/��h,��\������'���VR�Q{/��Z�IJ��Ms��;.��^�)ǋ�>���c����g��]5�ʯ��L�c�U�>�j��iv<P)��_;QW�n�?�պ��n���%G�I׾���r�iK i�����}/VR���C%�:s/����x��1g	������ôiK�h�/�����oJ����)�X�9:u�{u-v��pF�s�{Ea�7Ocٚ�9>��M������]y�8a0��#L�hʱ�o����NOQ'o��.�����S�z&P�~�2]���l}��F>��,��:��S�W�7�U���u�V�@{!l������_6C�+z��<�V�UⰧVR���h��ܫJ�B��ˏ4�q���|0�m�aȾ�ݦY�Ǆ��)��~sNȸk�(s�Yu���+���z,�]���|8m5K{�H��Z+j<C��9���n���{<M�X��>���Ǭ�W?)in��]���&�w�'G�e��äx���;�rb���!;�,�{=l����}�@�\�IW7�}��㇬�����F�����SҿL?�n�5uַG���uu]mZb��.M�9��T�zj�f'9�^4����B���P�/��x�����I���n�@ �Ǒ N�2�3iM�]}��l�UM�*q�Bڇ��ENF�:�{��o[�-m�j�j�~D��l�fzJ ��鋧~�+Z"���wv����w��j�7�#� :�~�a�Ah��i����D�+n^��Cw�Y֩�����u���xmh��[�D�o_�ft��H����J��P�X�D���!�~;����Ry��{����M���ڔ����'��G<�Y%�?nlZsm�Z�'�\�j���{�Тڏg��Ҏ���W�?nM��ˇ���yn��6U�vEF�B����^���T��?*�>ǣ�&Ls��D��ģ��'��`j2���g�j-N��u�z�\^l��+�0Jk�����n���k&���7����T>/����k�e�m,k��*�a\�^�w�~��yo�%�Fn�K��{��e�<N�%��O�V4��n?�\e�d����P�=��6i�>��,ǔ���#���~>��{�ޕS�#�G�G�)sJiM�m�վ�����ΩՁ�Z7�Y]i|?��v���}oXaY�9y��O���u�7�m%"9�G�����<��ϧ�N+��t�MN,ʌ������_��#n<��l��N1�l�ٱ=p��*OK.�8I�y�$U#��N�<�ױf�i��*��oy\�5M�s	�~<]�){\�t�S�C5�uO�U����㭀���C�yJ���������A�+�ۄ��=,�_�r8e�v����q��Z��o�y��V���r$wqװ�j�q�'��,�\T�I��\X�l�|Fv���ւ�L��.���z�Zb�r�Q
ơ�g�m��nX���9�r����m�����+�]
U�t��xS!�v���y�g5/*��ٟI��yɹ�|܇zi,+�'V��q�}�e�Pv��f,����,��`�Sj�m����;>7�~c���MYⷹM��~�(��z�������s����S��j{P`e�ʛ��)G���0��=\I����"~3�n<b݌�3�L�tL�*	��T��������z��\]W�<�(�����^�������?�:���xH�P�u�T�V�*�oK6��T`#u���̭�:�m���h�]9�X�aE:/q��F�grL-��4яK����'X~�����䕯�+$j�~�<PV`S�z�巀߀�E��N�\�a�g{&I�_�ϻWǗxui�L��g��Jq0S����l�!*+<9D�UK#�B:pz�����}�v�ҿ�<�:�3�c����"��e��p������_Yx���XK߮�����g��iK�?����Z1<��[uQz����Α�ŏ�kK��iO/W���ݷhI��v��gf+7�T�d@��	�~��4oQp�e����E�n��Gm�U�X��Y������d=m���✞�V"�QV���νg]@X���Uz��Zr�)[��)�ȁ�h�f�C��.-�m߼8Y�k΃K_%�ww�"�'�~�p�d��C"�b��зCw����*��/b���w�Y6�����V�S�g�X�0�حԾ�*w�����W��H<U�#��wa�;C�`����s9�F_C��za�����n�O�}�p�V.�Ӕ(�T�YwC�?1�E��oV���9��+Q��48LZ0q�	��֓�U���#�G]w����*�׾G&X"���󔉏Q�0h�Y��S8�A:����TT�ٷ��<x���C�o�o=�}��C5�SQ��9P��=	��*_�<;r���˸�����j�+àw>��+�vh�?V��Sn�>���<�\0��9����u��EI��}=^�=�cѣ��︝y�?٢|��`���w%lҤ��N�����,�A
۵$n�݌��94�-qx�S5�p�BՂ�\��&���W�`�Ȗ�m\���zk�M��O����}�D���o���Q\wZ#�];'��8��p������V0�z��{U�Ò���
F<Vڻ��m�݋_*'2߯#�1WB	�%_䵙��׾DX��>vŻ%w����q.�J�Ej<6@��y㺮*˛~���^�#�x��-凛�{�3Ft�ɒ]�^.�崙V�e�IR:Ń�Ld�:<�j�ߦ��r�U7�!�պ�J�asS�q��7��?�xb���Dq������o?����݂�'ory��܊�6r�I�%k4ɍ�D�x�MA~��������_a��d���ݝ9��5�򫬞��c�����t��^�Ԏy۵�ڪ�:���H�Մzm����5]r�C�X����|]X����;<��>+������ɟ�*����Z��Y@kJP?2x����Y��2�����,J:�� �:��?�t`*-��Ӕl]�azG�`[��K�&M���t��X����O��͡��ބ��=J��_rM���FUKb�N-���?�T�`?YW���)p1Xb�?c�ܟ3,���g������W�NW�j�M��'�.^f*(�w^�?���XU���k~�)�o-�ǎ��1,O��1�ʛ"�b���c2�Q:[r�{�h��_�"+�}Mјؘq&Mc��-�a�kQ��N�[���bsE*��o'������|֦�=Uje��S��8�����his����֕�W*J�
�jj�z�~��d�%t�6���EG7`�<���&�.��bYLx2g�{ұ]�:��/������7)P~25�Y��u�����I�������;�gH�z4���"~�s���?�jv>��#��G���n4m�xt��������\�+ϥ�9O�~�kH��>��ٴ���O�5��怟Ϲ�Jκ�C��E�(o��mO�p�b����V�<q����?�����F�%��.�U{6�-j��{�r�M��VEo��{���-k�)ɿ<����[>s��T����x}x��B�BE��&����oW����\-���l�C�j�{�0�],{Q�&���%\�Z	�d�Hϕ6�n'�難�MJ��!R�/ރj\ZgI���.�s����s�m#+�O��7~�i9��c���h�/�d�E�CԆ�^D���N��i�ɋ��8�~��7����\W���7�\��b<�Xy��
N�v����מ3�A�u>�Z�ɣ
�����)0��,=h/ꜻ㜤�ܛ��~��-���:H�a���1�[L9��;����pFzK�c�=���J~S'��q��b\�M>Ƿi_i��&��^���R��� �*��yi��F��Ãu��i#6�Y�����l�=�frTQ��;�\�!x�/`��'�؉;?�o����F2��W�f���d}߅�;���&u�|J��RL��'�|���N�k�kT�H��5V�B��o���{b���k�+� ]Wqo._q�<�ڻ��Zb�O^72��S�-B�^h��3aRV�|u����ʊAOxP��S�4y��b�L�"�l����e��#�w�f�O��xq����hJ���I��}�o���]�� 	�D?���s�;�OZ<L�~�W����+�A�ІҪ���v\[���=��4�Kw�i\>Ns�o��yi�k.@ӺO��0�F��=�t�E���Bs��q��OMmi:Z/�ۥ��g��k��S�_L4�|�L^��k<�"��r0�͡����$�P����H�.��&����x����J��-YS�}�m�5.U�K�	Y2�D���K���/�W<�������o��
��{gB|�$I<�?Ё�S�3��[����Q�ɱ<����]�k!�1s�c׮)�u��x|&���&�u�V��s3�&6��L�5�q���#�f�ՉG;"�]�w�T���M�q٘�>�w�H��k���]wr����CVO�>~>����.��K{�2��X�����N�>��n{Ɔ����r�Ǹ{z�a�4:���*	���)��&��&��Ð������h���Ӌ����R����oL��?����1-WC��rW`�O�Fs-��7׾�<�H����r���8�|N6��vO[ p
(䍄�K�pD�*��;�n���\������3�vefO��n*�����蚉$�49v�t�d�c���Ѻ����[��������<xpN7�X�/V���[(C#T��ڏ�n���L��е��Ѱ�\!�R�B瘽v�l�&�����w�Z1���Jo����菻����%��_�'E��S��	����[��(�*�V��5g�IP���y��&/��W��)�n;���e�o����m�"5_$T_K�?�k��wd�½w�^��;v�����.<Z��Y����M�+��l&q��K?a{7�kR��:����Y��1�I�B��W�_�헒W����Lm;3�>f��n���wK}���KJl���Y���)[��OM���s�2����ύ9%p�����s1�s�0+WVVn��e#V��8�K�Ju�Q�}뽂�jw.[,��>�l�΋!�:&����ȏ��fq�CAwf5?�$��شcC�≟��޶`o'�:��6�����P��/���h,&�Z �5��K�h���xʌ�]�񂥼��o��<{*���JF�A���鈸3R��0���0F9��fDzi����T��1mo�,E�*�B����b�^Y�n��D����{�`�8��'��cq�R�)9!�ܴ��/���T,�����Qj����q�z��1J:���ȋ�M��Kz�J��MZF�b����J-5�?�M�3#E�1��<������SW���ˬ��W�Ͻ:\5�9�����k�W�t���f���kxTv}Kh
���1��������1�|sB�U��I	�ʋ[�4e��܍����ȍ������,��ӵ�J����X��0 �Pvq��阃���ƈ["zx���s��n�\�y�']u���P��I�q��;����L�(����ٙNK�C;צ�S���\*�x��ZX�����R����������$N�+���M9�k=���x�'�w3Ft
���Y�Z�ex���:�E��F3o7Dϵ�0�Aܥ�����I�z��_?��1ʞ����.�+��.⣅.�)�N�n+#.n�k�,�@㾯�όj��PFTdh��0������e���u�bo�3ք���u�1b�GtX�i��e!ACؠkP��H8k���� 
y}xb]����`���,��fj4���=u ~�#
�O���X^�P�d�F�.8_�{u�Y�������~��t��"�#SA��IvF����X�kӛ�����v�e���<�j�ؖ�(���1�4?�����Ώ}L�"�-��M�<�zW@67'n�}c»����)=��*iکup�x�:')�)�I��3Η�J�	���a���%*-#�5|u����K���
�,�.�Fë���;�0킮o5n�c������|d���=˓t�!��?��|4=��d5T�n�ƺ��V���5oL�FFds��fh,t�Do�_`�;Kk~�2zk��,�s���H���&o���u�Ē���Z��0'4|^�)H#%-܊wBesٳgy; � CA{���i�&�[�b��@�'��s���כ��|��=���ҏ�<e� V�ЧI���;���ٟ���t�3��$��J����l��n��j�0+��^ʈQ�>�2t+��$�J�#��CW��s_�� ��D!_����=J��Ҁܺ�+4�Fޙ��@�J0$ѫI_�)8�X[#���Ǩ��}1 }��d�p#�h�ff��s�}��I�*$��e�c�SO%7m�����l01N2A������涊m�sb�aa�D$����ey�?�4yH���N���?{�0�rDo��I0�m�vo�Լ�*���(���g��Q�#��W���܇�z�]�4��M��
�@|]��1�O�����ِ�جB�;0��L����HK�8k4�a6dh�� ��Ak�� |������ȳF�T�'�����Sv�����ќ�h*��]��Dl�m X��/	����k�1�ȁ�Fx���#�ťqi��q8C�hߧƤ\��^}*|q��D!#�?߇r�ء�ɇ�Ih5�۫��uS���т�U����az�BQ5T��S�6��o&!���?��x���>�9彣�Y]@>:��1iD*��Ԇ*;B� ^��E@o����s��t@+���=Ϫy�c�V�mձ
�a�ֆ���lH&nw�sr"GtΜ�����0�fD�q���X��vd@AJ�s���Bt��S�mD��[��*}O����e^����~d�� ��@|"bEY)��Wֻ����YnS*����|`1e���|r��z�6R���lj�W���8�Z��~���������X�s�<�{��:�p'����Ǆ|9�5�8�(�R��hG��?�^>�n�K@��{���G��� ~�T��+��)`�"Gr.�aj{�Ėd�i?}YiF4��:�}�ⶣ��!�[�f�}o�P(j�[oޜl��P(�P�3z�=�`ɢ	r2�]3��s�#Q1����\wv'JR��l{� f�Y	���b��/��O���wļ��j-�߳�l���٪3�@h�V��!�#橭V�>�Ě�}����=��6�Iy��ȉLZT�b�w�	A�ڣ��Î�x�IpP{,.�(����v&�=|8�-����X��J5=�퉡��6�n>�����5�ak��ຄFF��ng�=�����Mǭ�'��O%��)`��ec��|V��#�'I�b/�x��񷿞�'���D�"L��{{�'����lD�3����S�<vsߍ*�j��ԓu���(��ܩz��+U�C�?��P����폸u��G�޳]�JBv��H=8.����}�����S�A��9l>�D�<�w\-�t�#K���������"#��S\G��Z���=�u�d�r~lpI�����G�aO{��ͽ O���B	c���@��o�a�d�#��j��3f����}tƿ>vcVaVaVaVaVaVaVaVaVaVaVaVaVaVaVaV��z�?
����/V��V�.ۯ"1�A���^�;, ��w��k���:�ή���:�ή���:�ή���:�ή���:�ή�+Zw6D��(��t�|��~�vv�]g��uv�]g��uv�]�/\n���׻ �_�2�ή���:�ή���:�ή��6g^����\P�g�gbE�3驖I�Yh�&��-iJ�W�������*�MƼFtc�=v?�u��k����_���j}�bh����z�Mm|����l�g��+��mg��50k`����Y�f��50k`����Y��_P&ߘ��d���7���|K�<��-���(/'��v7���2:������wb�wI���|/����r�yc�
s0ڈ����	O�w:�������ʊɦ|^orDor���?���B���RxE|�]�,9�:1y���C�)F��0�ɸ��?��/��,��9o�FM��:i����i���~T��b�\#�{OﱱŒ%�e��'*����0�'>\ՈY)G=��-�H�X���I�*�������3T�W�| _��WQ�ĤFA��x�~�DRY����NL����jIc�b�Z؇�T���Pu�z�&����X��HN�b��е̠"dF�,*��r	>�� T�w���pib9��nvb��ɸ�_Ȱ2�����&����߅?oUC�,E�0����y��|�퉊
�󏼃%��Ɵ>��iQ�rE_��(h�ہ}����)�7���|P�F���`&Lp�rl6t�P;'I(���=�`�E%��~�O�����{)�X�](_�F��f���N�r��\��kޝ;1y'׼���2J�؜��ڠF�ܪ���&�a�np1�/ӡ�1"�
�n���'�Q��Ȱ�,M��l���Tx�(�����%��>���?�SL�u�eQ=g,�∽���qΑ��Q.��!���TB����.��$����'S��R@ċ�	�G�$� e�B��(���Xi��sl��w�nF HB��y3ԑY6�}9��t�O����g��%N�* Ჷ�s��n��#��+�3�#_~���>�3 F�#n�Cʼ��<�����]�[�!�`�𶙡0����%`�O�y�ϟ�d(#�5�9|r�)�3S�?��Kt�Iq���nHQ�*��ݽ	�������8TN37�D�!t�7����l���q��p��~Ri�yG9��Cԝ�I��2'�*(�Q������F�, "r��Vt^)�/���-�����QVe�ڂ���D��%ePbMr�T�2�&
/���$�d�Ex5�����L5z�ո�����Y���Ah���f(��iAI�1�t��oj�ā����/�d��#da�'Ya9C���`)�K'�Ā�5�#�QR�/��30
���L��ڸ��tP ��Ӝ�IBT(��)(���q��t\���ÖL�I����� D?�J5�K'�.�U>1�d��Qo\�+(�DdREPܷ�<Ce��U����� e�T�V� �ԮAҍ֙��.�+C�T���Du�#���w��2��əR�t�֔���݊	zc"lT�:�����b2Ȭ�����>��C��6�s��U �Np3�u�L���Qg')�ŏs����nO�Q ,�`41�H�5� "�5�Te�L���	FʕO'&?ч�>�\+} ���F�L-��"����F�́�-�ٱA�]��WPg�D�VC������98�﬎�B�Q����3G�w�,)Q;<4�ϟ��������IK�0lx�>s�l���������N��V&��57���!��&(7��L��upX�ߐ��d����q� ��>SC�zh��w�ߊ�0�3�^�A㜭35i��12��*]?�,7�����wa�S� q�Iy�3A�v^E�P�2m�;ᝉ3ѐ�
L��͠�z�D1p�DA_Tğ�NVf�Pј��)���qj?�r+���(Cqa?�\�.=�u�M8Ȕ����	���<�F?�PCE��qxp�L+�Mx���H�S*d$�q��������d�<.�a������o\
�#�`ɝ���qѡt����X3tdt�#�6@GF�؄7�#>�
N��J��������ѱ	�0i�DV��Б�R�<�����	�+�^�A;�� :��������ꭔ�V���̡k��Z�2����׆f�<8�C�����:�Q��@����q���KG�A�Aߔ=�L�+��S
�����F��[��鈎�@��}))�a������l�����«7�5���u�'�53t����Eo��a��T*}�����I�����|Vv;x�`�8������h�S�+g~P��4t�I-U��wH#g��ۣTj];Q��\D�}x9�H0��; mF[d���[r��	� �g� �� �_��'����n��4���.�1���H#_[Qa�1��G�Ժ���]zR!�E���O��U����Ol�~�K%B� �Q�����2�5h��-e	[�bOQ�����|�O��>�Z�'BI)·r8n�ՙe��4�_6T��Q���&�9�}����� ��^8&o�N3�������'P����g\���`hC%�}��%P�i3���@Q�l�5�m@ABܘ�����م�l�ɏT��Yd�@����cXLPv�#��CVW�2����d�eP��N�����f��pP�gtȍ�ƕ�����������"��YܸG?��ɹ��?C�S!��wg����J�C��-�h�5�!��yS*���U���ȡ�D����C>�T&���^- �&�V�7���'Ɠ����H	���ߐ�^�E>5¬5�v|�BD	Qb$n������/�|�Ռ��F�r�u'����\���F�y���7/����F�\�An�z����qo|*���$���+�9���������36;�ȫ���p�re_���:~R��D_������v�Ers*g�s����G�f��L�N�HS�D���wKQ�%�@���Ar`���ޕ��Gy�����r.�.B%��3ݐ��?�a?@�o�HmӝI%�t��oVָG��S��:@u���%�� �����$�c&MG����Q������g�~�x��b��"u����
 �9�34�T�r	�����3I߹&��1��b{��w�@��T�u�f��c��ȑ WVQ��19�}���)���:�|~/��;�zO,p�#����b$��޻�=`���zo�z������`��*��,���\4�^9�Q�G��Y�ȋ��1ȡ7�c�ģ�NTQ��,�s'�5h�(TU/�@(��J�	0灛{�I'~��M0|&+y�����>�N���O� ��0��Kj~W��$a�'�L�K;QY.���Uǰt�O �*��~ �W���Z��_3�F��@�x� Jsа8���%�Tu A�Y���p�ͽ�d�!���2Q6�}��d!��O�42@X"��M턽J ��d���s_S�׊��A(�(.�*�^&C6CR,�2l	#MG(]�@2_$�F�ޢA�Yr�0���.i� 4<��R�W�$�E�!+]ڎD_A�;�u��Y��h;��N2��:��]����J��!K����-c���"�!��%%�ˬ�;�ډ�o�{õG3$;2(�U�b?��$F�#�E*]r��fGجQ������߲�BBpݡ�f�:K�&� slD}3W�N�z+~�D~H����K��sI	��^���.)��ώNm�{��=��܈z����F!�A+�Cw*���fT^�p�3�	z%~|�	y���M�#ݸ�tIl+��c�� s����(�q����-�� �����qX'p�n�鉁��>�I؋d�H���2�e3���Jګ{=X-�[zs��Q���Y{AF�A�*�1��L؋���n{�,��{�\��ڤR/s=�HF2M$�YiSK6��#���{7�#{����"�˼{Af����D����Z���)G�"^����\�'��?��"������b��(�%��rȗA	!�B���U��2�f������-FSR3�w��@0#u&��9��߼�$6z��KfX
��RtĎu�&"�:��f�����tC��9�̇�v�._���X	-Qף;@�r'w�є�:Rż�Ԥ��"�	|9V(ƕ�(@��^��IG�a����8���蠨��h�$�1m!����=�����A,�B"D��Y,�l��� �1��/!�_���5��)���|��Y(ʖ����I�e������)�/q���;m���QO2�iY^�EV���r醌�`�����dt�T4���yg?�_��9�~��~k۝Qhs�P��Y�12Y�2w����b�e�a81;�)R�@syM�q0����G"� t�����5�B�`��cq�d3:j/�ƚj?B>4�e��C(��HbO�RC�E$��˭�' v��-*4,��"�hX�Pǰ�)u!��Fj�j;r��5h��f�Є�(C;Cmr���iY~oL0h�\I�����a=8}M�VDZ��Nk;�p�7�S���BC��Z������s�[�B�nPAִ��Kj�3=/���N��9��(�Ks �	���0I,�-u�Hڔ"��8@j������1@�����~b�0��Ajw�!���?>�f� ;��\N�I��H��U&��&�r���ć�*b�~�Xp���A8P����zp� ^,��	�p»Cd��^��l�����^���_��K��[�����(�}/�H#��؉~œ���!�~^*�sA��S��,h��\W"��,-��q�A}��Wd�w7��a3�ڋ׼$W��ari���� �]�"]��L���D��כX{H)��:N�"�.�T�;,sp
�&�#}j��R�Mkp���a/��Z�S�	8�pk�AMw
HW�2G�i8ő�5@J��"�ӹ�S@*����zrZ��7t�HqeM�c�^й(����C��q-CK�h��ʐ��A�l
~[��&4�cI��V�HQ2��6��؂�]d�w�.�V�܏��7�2ut�?��&n�e0���2�g|�B2%\c�[-#�B�3���yK���c���{�'��)�Ռ>؋dx�wܪ������\�^�7�} z�^3<��2�g~�B2�P�!e& W�h���$;���>f�}z�p=�!B�W`/��ؚa�2�fx�^Hw�M�w��e��^8Z*O�L�5��=��C�$��8��[K�z����G��K���83c_�l,A� �%���6���"��4���1hkt�}�YZ*�*��V�F,��%\Y�}�PH.idN&ƪj��&Q���Z>���A���~[ɕEe���s�K�, �����$�md�Ҙ�AÑ��Mn�NɅ�N�#�c��M��c������O����K"�2n�\ko2�[@�����������<#�!	�w��&A���B��&h�� ������jЂ�W��(m���DH!���@�f��3\�fn�� ��e˸�P'�=^� �N�8IL'�j{�n���B�A(�^�s��'!��pԗx���9u���{F��qV��X�c_���I�J��C,p����]�2��B%�b%Jˉ��:�-�F��������z���<Y繲Rz���	���1(R�~��bh�3zWAoٍ~0\���bYxy�37G@�&�b�߁�*
��r���pG�.�sWֳ�����y?��k�O�E��`?�w���rsą���%�2D�I�X
QO���|�C}���M5s*ʅ˭u0�|-�:�0R���ڶ:!�C}%I�R��\��-�6�ؑ^�+��g�Ok3K���:�D�#�B3��Ϲw�Y���y� �t���[��[qcB$��>f��������^�'ޮOQ_��<Q�80�E�o��Zd�+�<�́1�Hx®#�����a	0�+��a>ai-��E�p���a^�e��~^�m��0{ �2R���f��L�$���90!�Wq�4�V�K*��i�8�S���B�r��0�?�������p��'s:��ӾB�T%吡VѨ�-Λ�SH���:$��>�"�
�>������,�H"p�2��V�3��(R�/�G,����A2�~�xH�w����J�*��'���~��$����%��`j�^����
IR��]���� Yx�O`8d0�,��Ӛ���u��Fh8����\�k���[���Dϣ��W����-�㋨[�}�+Ε=_���D&Ae�!��	�P<!�'!<<�����܈��U{�m%����֒�� d8�_����|(��3�6E��[�Z;�3�Ǡ��!�>g8�{�nPc�!��N�A�((E)�f��j�sGw��!T�<<H�Kkĉ^uB��7�-u� ��Kg}QvE��f���X|�s�(�-<���_ο�w��";(�Γ:���҂���M��e~�/�
��{������J�Q���:g�l�5h-P��xi輦~��F��f���,��#^����rYZ^��يF�<nP�+;N�E�\��"���@��A��=UÀ�[e��F�z�3�B�mB 4�`@�g�A�N|C�*���ĩ8��,-s��-�K��{��b���rnD4%�4��@0��|�^��ږ(��
-nY�,�3q��XZ�H��e~ځ��f!W�g-#�>
�p=5�{E���-�ӎ�e�Ұ��~��g\O��'9� �����_-|/t�F���[8�p�p��,������O�$�U�����ވ��0x8�F�t���ކ��^gY���kv��/�!��B�����Ӗ�v�[H��Ar�vnD�h�!E���E�#B�=K+E��y����zrT����<�^g�ۜ��M� �G�F#���FYێ����Hb!}Ή]ڡ��tfs�3��K����D�Q��J�ڐ��(,�@JG_9�r��"r6j������@�1�"� ����#ކA�)�PGצٲ�e$���XQ��+��b�E��r[�sO��9��>�=�yϹ�f�n��R���:f���g�A8�3����Ƨw���s#$3B�N�_���Ƭҹ+�O�W���@<��� �2�* &�u���UR�w˅��Ư��B��)"�I?%��g��{͊��y�sʂy�CB׬�OȲv�ID��c�aD�����R�O\Ԥb���W�6�����S�^���g�z�=���E�B�7�j���a^�R���0p���M�WlQV��*�K�?o�>��{��^�g�
Y�Z?����9g��Ա ����-ɏLH1��A�WZ]n�M�8�=�]��0h��Xh\��
��3|D@n�o���u)�jd�i�������R�O�!��t����Ъc!j���'�-�x�ʜ?z�ڏ�46;��|<�������p��;tE��p���t���f�_����nu̖���+��u�ަ�cs����z���9���T�0�V����<g;b��V[Ƹ|Y��6�a��QY�$��x Qev-m4�h�,�@�q����S7!5��g-�7�h���̸���dÌ�cxo���`��|�]K�R����º��g�
l��3<�+�Sf2+bhU�Q�4�zݤ��+�_��u��Z���R�a\1H�����"RC��~	�R����ٰ\������^O�&$+n� �Ld�b\�,\ i��)5�J_����ŤtJM����f����P�{�\o�R2t#�e��ܪӆ��\y�a��];9��g�PK    {�XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK    {�Xt��  �%     jsons/user_defined.json��N�H�_%�4Ү���~� =�H4�͎4B�����`���Q��4/�ϴ�N���4̎vE��/�_�*��:�����2&{I����!fyC2M>�j����)N	\Yծi�J�~�zsrb��gg��w��0"��������@�dlV��:���=n;���b�I����D9��� "w4D��΀ø�U�\o����.�pn��Bb�$�qm	r3Dc���1��e��[��Q����פ����ra��a�R�|��ݭ���oo��f6�"�T��Q����aښ�*o�|�/����'��J�Y�?�<�쭫�da]l��rr�|�����8yT};�7����iG�>U��� �v��������
^�7�T��X��+m�o��&|�SWˢqC���3���S0v�}����⠼Z�v���E���"�^�⧺��f�C�٢ά_�U�����'GE��g�������x,�Zy%-b��+�!-�B�xh�$���c=�S�X_��I@��~��%P�!b��߽�c���Z�:/��������}U�U�\,`vKYp�VJ��YLҎ�%�t,��Ac�� �� -�_E=��[���5
v3�=��ګ����IEǔ<a�����}�~��I��~�L�����	�1J�,��zP�ue�(Y���AU�UU�TŰ��j�Q��"�슚g��n|ţD/�ڐ���Q�3<�i��<�$���Ŋ����BE�y������q�?�â]��8ן�a�.O��)}<O���U{��#egò=L�q��]�t�"t��εV,������e��� О�%��CK{��+;_hO�R#eͰjO��#U��j��6j�QUê]�(�*�U����`��p��=y��T��'q��xў�%F���zr��:�I^j�*���
/��Q���3�!Ǵ���˨�>0vS`�Hi6k�A)���lS�LE���|i��\�y�/&o�|�X<��bUVʭ�mV�wF���H�9c<��(#P�f�Qu�τaTe�:����(i�,��̎�1�;#���I�O��7)�B�i�Ri�k�vat��o�/�v�Ęg,	�YK<����/O(�������8�D)����s�J�@�TQֆ���nZc���i��&���	"�����z���/�}$��54H��]�in2��9��/�}t��por~]N�uM��%.���wD�6�y�QX(H���HeV"b�@RDC�S��� :���e=�k|/�F3�C�o&��4Uac�f
�Dt�ڣj�����=�4ժa�n4a��CRXu>�Y��X��3���B�#�1�Ѱ5��Ek��g#-%\��=qs�|��U��6N�������;�������pyiX	��� 9E<X�Uc$8�e�ς���EUk��%	� kx���
�3�����Z��F!�3@C���d���s�x�+�������@��u����	X���CJ�A"@�"�<�sX:�r�����Ra߮����_K��D�Z�0����E��$�vlM`%��@���f�I&�73X>�H�vx}p?RD�ͪY�@���(F�r
���~�t�)�[�Q0��#�'y������pl���rj�co�������} �'�pf���ox��H|���	�uq��y����~�����5F'8��%��Ϳ��=������8z���k�I}�b59�&���;�����Q}݋�yM��f7% 7�r�,c�`E���5"�F�׈�^ "\~�PK
    {�X�l�@  �                   cirkitFile.jsonPK
    {�X��U
a6  \6  /             m  images/0287c76a-3da1-471f-86e7-79c7d2df61ef.pngPK
    {�Xyɜ��  �  /             H  images/110f4c69-ce42-4daf-8800-65b9db14e3fe.pngPK
    {�X�䓶� � /             �d  images/132fbcdf-34e4-44dc-827d-09a965026955.pngPK
    {�X�?HU!  B#  /              images/585092fd-6de4-462f-8499-92296fb2c536.pngPK
    {�Xd��  �   /             �: images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
    {�X	��#u } /             �Z images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
    {�X��Xc_@ �d /             )� images/a9ae5602-6322-48a1-b803-2efd75c9b3bb.pngPK
    {�X+L$��� �� /             � images/aad47697-5cf4-402f-a095-abba84463b41.pngPK
    {�X����<  �  /             ��	 images/bdd7c0cc-86d6-4eb9-abef-3fcf444ec41a.pngPK
    {�X$7h�!  �!  /             �
 images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
    {�XXs�銙 � /             �#
 images/cf59327f-2b20-4f20-97ad-1ec426c5b43a.pngPK
    {�XP��/�  ǽ  /             �� images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
    {�Xt��  �%               �o jsons/user_defined.jsonPK      �  w   